module tb;
parameter data_w=8;
parameter C=12;
parameter R=24;
parameter D=24;
reg [C*R*data_w-1:0] m;
reg [R*D*data_w-1:0] l;
wire [R*D-1:0] s;
reg clk, rst;
wire [1:0] status;

ldpc_core #(.C(C), .R(R), .D(D), .data_w(data_w)) X (1'b1,clk,rst,l,m,s,status);

//A set of test data
//WiMax 1/2 rate,576 bits encoded random data

initial begin
	m={8'd0,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd7,8'd26,-8'd1,-8'd1,-8'd1,8'd41,-8'd1,8'd66,-8'd1,-8'd1,-8'd1,-8'd1,8'd43,8'd0,8'd0,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd49,8'd39,-8'd1,-8'd1,-8'd1,-8'd1,8'd65,8'd7,-8'd1,-8'd1,-8'd1,8'd0,8'd0,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd72,8'd70,-8'd1,-8'd1,8'd59,-8'd1,8'd94,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd0,8'd0,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd51,-8'd1,-8'd1,-8'd1,8'd43,-8'd1,8'd24,8'd83,-8'd1,-8'd1,-8'd1,8'd12,-8'd1,-8'd1,-8'd1,8'd0,8'd0,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd47,-8'd1,-8'd1,8'd2,-8'd1,-8'd1,-8'd1,8'd73,8'd11,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd0,8'd0,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd18,8'd14,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd53,8'd95,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd0,8'd0,-8'd1,-8'd1,-8'd1,-8'd1,8'd0,8'd79,-8'd1,-8'd1,-8'd1,8'd82,-8'd1,8'd40,8'd46,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd0,8'd0,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd72,8'd41,-8'd1,-8'd1,8'd84,-8'd1,-8'd1,-8'd1,8'd39,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd0,8'd0,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd25,8'd65,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd47,-8'd1,8'd61,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd0,8'd0,-8'd1,-8'd1,8'd0,-8'd1,-8'd1,-8'd1,8'd33,-8'd1,8'd81,8'd22,8'd24,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd0,8'd0,-8'd1,8'd12,-8'd1,-8'd1,-8'd1,8'd9,8'd79,8'd22,-8'd1,-8'd1,-8'd1,8'd27,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd0,8'd7,-8'd1,-8'd1,8'd83,8'd55,-8'd1,-8'd1,-8'd1,-8'd1,-8'd1,8'd73,8'd94,-8'd1};
	l={-8'd20,-8'd5,8'd28,-8'd72,8'd42,-8'd33,8'd48,-8'd44,8'd29,8'd11,8'd74,8'd12,-8'd36,8'd28,8'd6,8'd87,8'd20,8'd32,8'd3,-8'd63,-8'd32,8'd2,8'd31,8'd5,8'd28,8'd14,8'd17,-8'd33,8'd23,8'd5,8'd17,8'd2,8'd42,-8'd6,-8'd26,-8'd49,8'd56,8'd31,8'd27,-8'd17,8'd43,-8'd29,8'd20,-8'd60,-8'd22,8'd20,8'd27,-8'd16,-8'd4,8'd8,8'd42,-8'd27,8'd26,-8'd6,-8'd4,8'd27,-8'd36,-8'd35,8'd46,-8'd20,-8'd34,8'd25,-8'd34,8'd3,-8'd6,-8'd44,-8'd36,-8'd37,-8'd18,-8'd10,-8'd23,-8'd51,8'd36,8'd21,8'd41,-8'd23,8'd13,8'd39,8'd8,-8'd11,-8'd58,8'd22,-8'd7,8'd6,8'd42,-8'd70,-8'd30,-8'd38,8'd11,8'd11,8'd15,8'd10,-8'd25,8'd19,-8'd30,8'd32,-8'd13,-8'd40,-8'd20,-8'd34,-8'd42,8'd46,8'd1,-8'd1,-8'd9,-8'd60,8'd9,8'd42,-8'd43,8'd48,8'd53,-8'd4,-8'd22,8'd30,8'd48,-8'd48,8'd27,-8'd26,8'd35,8'd32,8'd3,-8'd55,8'd7,-8'd15,8'd16,8'd6,8'd1,8'd12,-8'd57,8'd23,8'd34,8'd9,-8'd10,-8'd73,-8'd18,8'd35,8'd10,8'd1,-8'd33,-8'd28,8'd50,-8'd4,-8'd18,8'd14,8'd29,8'd39,-8'd19,-8'd24,8'd23,-8'd23,8'd57,8'd15,-8'd47,-8'd1,8'd26,8'd23,-8'd24,-8'd11,-8'd31,-8'd8,8'd55,-8'd5,-8'd62,-8'd26,-8'd62,8'd39,-8'd17,-8'd56,8'd29,8'd10,-8'd33,8'd10,8'd14,8'd13,8'd28,-8'd19,-8'd21,-8'd22,-8'd27,8'd0,8'd51,-8'd44,8'd5,8'd4,-8'd49,-8'd44,-8'd6,8'd45,8'd13,8'd51,8'd22,8'd6,8'd24,-8'd3,8'd46,-8'd11,8'd45,-8'd39,-8'd13,8'd58,8'd1,-8'd19,-8'd51,8'd44,8'd34,8'd46,-8'd14,-8'd37,8'd10,8'd62,-8'd26,8'd15,-8'd38,-8'd45,8'd15,-8'd10,8'd28,-8'd30,-8'd4,8'd42,-8'd52,-8'd67,8'd46,-8'd65,8'd1,8'd11,8'd10,8'd38,8'd77,8'd25,8'd9,-8'd31,-8'd30,8'd47,8'd39,-8'd14,-8'd15,8'd35,-8'd23,8'd11,8'd22,8'd31,-8'd20,-8'd14,-8'd16,-8'd66,-8'd1,8'd35,8'd18,8'd15,8'd28,-8'd25,8'd2,-8'd29,-8'd39,-8'd4,8'd35,-8'd76,-8'd37,8'd4,8'd22,8'd25,-8'd16,-8'd49,8'd0,-8'd15,8'd1,-8'd14,-8'd55,8'd44,-8'd41,-8'd36,-8'd35,-8'd38,8'd22,8'd20,-8'd17,-8'd33,-8'd22,8'd23,8'd45,8'd50,-8'd11,-8'd17,8'd31,8'd22,-8'd21,8'd39,8'd11,-8'd47,8'd11,-8'd45,8'd18,-8'd56,-8'd12,-8'd46,-8'd30,8'd53,8'd51,8'd26,8'd26,8'd11,8'd1,-8'd21,8'd38,8'd37,-8'd37,-8'd20,8'd1,-8'd16,8'd18,-8'd6,8'd14,8'd55,-8'd22,-8'd25,-8'd47,8'd22,8'd43,-8'd30,8'd15,-8'd5,8'd4,8'd42,8'd12,8'd58,8'd47,-8'd45,-8'd48,-8'd13,8'd31,-8'd17,8'd10,8'd57,8'd16,-8'd37,8'd100,-8'd41,-8'd31,8'd69,-8'd11,-8'd29,8'd13,-8'd28,-8'd2,8'd61,8'd17,-8'd8,-8'd71,8'd1,-8'd41,-8'd7,-8'd34,8'd38,8'd61,-8'd22,8'd18,-8'd2,8'd5,-8'd5,8'd56,-8'd3,8'd43,8'd76,8'd5,-8'd28,8'd5,-8'd49,-8'd11,8'd24,-8'd3,-8'd5,8'd58,8'd2,8'd3,8'd18,-8'd45,8'd36,-8'd34,8'd15,-8'd29,-8'd32,-8'd35,-8'd32,8'd32,8'd27,8'd61,8'd9,8'd4,-8'd64,-8'd5,8'd52,8'd60,8'd29,8'd10,8'd58,-8'd37,8'd37,8'd47,8'd45,8'd35,-8'd22,8'd50,8'd6,8'd11,-8'd12,-8'd37,-8'd5,-8'd12,-8'd52,-8'd21,-8'd18,8'd35,-8'd6,-8'd60,8'd16,8'd13,-8'd31,-8'd20,-8'd47,-8'd16,-8'd11,-8'd15,-8'd38,8'd24,-8'd7,-8'd31,-8'd34,8'd44,-8'd12,8'd8,8'd21,-8'd33,8'd9,-8'd35,-8'd41,-8'd25,8'd28,8'd34,8'd24,8'd44,8'd25,-8'd11,-8'd7,-8'd28,-8'd1,8'd34,8'd29,-8'd21,-8'd18,-8'd13,-8'd20,8'd2,-8'd7,-8'd50,-8'd18,8'd43,8'd19,-8'd1,-8'd28,8'd12,-8'd42,-8'd15,8'd9,8'd25,-8'd51,-8'd39,-8'd21,8'd39,8'd37,-8'd15,-8'd27,-8'd4,-8'd42,-8'd45,-8'd30,-8'd17,-8'd18,8'd13,8'd14,8'd3,-8'd38,8'd36,8'd24,-8'd10,8'd32,-8'd11,8'd52,-8'd30,-8'd35,8'd39,-8'd34,8'd31,8'd55,-8'd31,-8'd19,-8'd3,-8'd8,-8'd32,-8'd66,8'd31,8'd11,8'd70,8'd20,-8'd28,-8'd5,8'd13,-8'd16,8'd11,-8'd25,-8'd2,8'd2,-8'd42,-8'd17,-8'd28,8'd3,-8'd24,8'd20,8'd29,-8'd45,8'd43,-8'd15,-8'd4,8'd63,8'd40,8'd30,-8'd7,-8'd35,-8'd1,8'd14,8'd26,-8'd51,-8'd29,8'd25,8'd0,8'd25,-8'd18,8'd16,-8'd22,-8'd35,8'd24,8'd14,8'd30,-8'd45,-8'd6,-8'd12,-8'd46,-8'd47,-8'd63,8'd7,-8'd37,8'd44,8'd29,-8'd24,8'd43,8'd12,-8'd5,-8'd17,8'd32,-8'd5,8'd15,8'd22,8'd16,-8'd18,-8'd17,-8'd29,-8'd1,8'd24,8'd59,-8'd62,-8'd6,8'd32,-8'd27,8'd72,-8'd19,-8'd1};

	clk = 0;
	#5 rst = 1;
	#10 rst = 0;
end

always
	#5 clk <= !clk;

always @(posedge status[0] or posedge status[1])
    #50 $finish;

endmodule

