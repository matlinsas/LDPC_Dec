module tb;
parameter data_w=12;
parameter C=12;
parameter R=24;
parameter D=24;
reg [C*R*data_w-1:0] m;
reg [R*D*data_w-1:0] l;
wire [R*D-1:0] s;
reg clk, rst;
wire [1:0] status;

top #(.C(C), .R(R), .D(D), .data_w(data_w)) X (clk,rst,l,m,s,status);

//A set of test data
//WiMax 1/2 rate,576 bits encoded random data

initial begin
	m={12'd0,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd7,12'd26,-12'd1,-12'd1,-12'd1,12'd41,-12'd1,12'd66,-12'd1,-12'd1,-12'd1,-12'd1,12'd43,12'd0,12'd0,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd49,12'd39,-12'd1,-12'd1,-12'd1,-12'd1,12'd65,12'd7,-12'd1,-12'd1,-12'd1,12'd0,12'd0,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd72,12'd70,-12'd1,-12'd1,12'd59,-12'd1,12'd94,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd0,12'd0,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd51,-12'd1,-12'd1,-12'd1,12'd43,-12'd1,12'd24,12'd83,-12'd1,-12'd1,-12'd1,12'd12,-12'd1,-12'd1,-12'd1,12'd0,12'd0,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd47,-12'd1,-12'd1,12'd2,-12'd1,-12'd1,-12'd1,12'd73,12'd11,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd0,12'd0,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd18,12'd14,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd53,12'd95,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd0,12'd0,-12'd1,-12'd1,-12'd1,-12'd1,12'd0,12'd79,-12'd1,-12'd1,-12'd1,12'd82,-12'd1,12'd40,12'd46,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd0,12'd0,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd72,12'd41,-12'd1,-12'd1,12'd84,-12'd1,-12'd1,-12'd1,12'd39,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd0,12'd0,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd25,12'd65,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd47,-12'd1,12'd61,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd0,12'd0,-12'd1,-12'd1,12'd0,-12'd1,-12'd1,-12'd1,12'd33,-12'd1,12'd81,12'd22,12'd24,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd0,12'd0,-12'd1,12'd12,-12'd1,-12'd1,-12'd1,12'd9,12'd79,12'd22,-12'd1,-12'd1,-12'd1,12'd27,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd0,12'd7,-12'd1,-12'd1,12'd83,12'd55,-12'd1,-12'd1,-12'd1,-12'd1,-12'd1,12'd73,12'd94,-12'd1};
	l={-12'd20,-12'd5,12'd28,-12'd72,12'd42,-12'd33,12'd48,-12'd44,12'd29,12'd11,12'd74,12'd12,-12'd36,12'd28,12'd6,12'd87,12'd20,12'd32,12'd3,-12'd63,-12'd32,12'd2,12'd31,12'd5,12'd28,12'd14,12'd17,-12'd33,12'd23,12'd5,12'd17,12'd2,12'd42,-12'd6,-12'd26,-12'd49,12'd56,12'd31,12'd27,-12'd17,12'd43,-12'd29,12'd20,-12'd60,-12'd22,12'd20,12'd27,-12'd16,-12'd4,12'd8,12'd42,-12'd27,12'd26,-12'd6,-12'd4,12'd27,-12'd36,-12'd35,12'd46,-12'd20,-12'd34,12'd25,-12'd34,12'd3,-12'd6,-12'd44,-12'd36,-12'd37,-12'd18,-12'd10,-12'd23,-12'd51,12'd36,12'd21,12'd41,-12'd23,12'd13,12'd39,12'd8,-12'd11,-12'd58,12'd22,-12'd7,12'd6,12'd42,-12'd70,-12'd30,-12'd38,12'd11,12'd11,12'd15,12'd10,-12'd25,12'd19,-12'd30,12'd32,-12'd13,-12'd40,-12'd20,-12'd34,-12'd42,12'd46,12'd1,-12'd1,-12'd9,-12'd60,12'd9,12'd42,-12'd43,12'd48,12'd53,-12'd4,-12'd22,12'd30,12'd48,-12'd48,12'd27,-12'd26,12'd35,12'd32,12'd3,-12'd55,12'd7,-12'd15,12'd16,12'd6,12'd1,12'd12,-12'd57,12'd23,12'd34,12'd9,-12'd10,-12'd73,-12'd18,12'd35,12'd10,12'd1,-12'd33,-12'd28,12'd50,-12'd4,-12'd18,12'd14,12'd29,12'd39,-12'd19,-12'd24,12'd23,-12'd23,12'd57,12'd15,-12'd47,-12'd1,12'd26,12'd23,-12'd24,-12'd11,-12'd31,-12'd8,12'd55,-12'd5,-12'd62,-12'd26,-12'd62,12'd39,-12'd17,-12'd56,12'd29,12'd10,-12'd33,12'd10,12'd14,12'd13,12'd28,-12'd19,-12'd21,-12'd22,-12'd27,12'd0,12'd51,-12'd44,12'd5,12'd4,-12'd49,-12'd44,-12'd6,12'd45,12'd13,12'd51,12'd22,12'd6,12'd24,-12'd3,12'd46,-12'd11,12'd45,-12'd39,-12'd13,12'd58,12'd1,-12'd19,-12'd51,12'd44,12'd34,12'd46,-12'd14,-12'd37,12'd10,12'd62,-12'd26,12'd15,-12'd38,-12'd45,12'd15,-12'd10,12'd28,-12'd30,-12'd4,12'd42,-12'd52,-12'd67,12'd46,-12'd65,12'd1,12'd11,12'd10,12'd38,12'd77,12'd25,12'd9,-12'd31,-12'd30,12'd47,12'd39,-12'd14,-12'd15,12'd35,-12'd23,12'd11,12'd22,12'd31,-12'd20,-12'd14,-12'd16,-12'd66,-12'd1,12'd35,12'd18,12'd15,12'd28,-12'd25,12'd2,-12'd29,-12'd39,-12'd4,12'd35,-12'd76,-12'd37,12'd4,12'd22,12'd25,-12'd16,-12'd49,12'd0,-12'd15,12'd1,-12'd14,-12'd55,12'd44,-12'd41,-12'd36,-12'd35,-12'd38,12'd22,12'd20,-12'd17,-12'd33,-12'd22,12'd23,12'd45,12'd50,-12'd11,-12'd17,12'd31,12'd22,-12'd21,12'd39,12'd11,-12'd47,12'd11,-12'd45,12'd18,-12'd56,-12'd12,-12'd46,-12'd30,12'd53,12'd51,12'd26,12'd26,12'd11,12'd1,-12'd21,12'd38,12'd37,-12'd37,-12'd20,12'd1,-12'd16,12'd18,-12'd6,12'd14,12'd55,-12'd22,-12'd25,-12'd47,12'd22,12'd43,-12'd30,12'd15,-12'd5,12'd4,12'd42,12'd12,12'd58,12'd47,-12'd45,-12'd48,-12'd13,12'd31,-12'd17,12'd10,12'd57,12'd16,-12'd37,12'd100,-12'd41,-12'd31,12'd69,-12'd11,-12'd29,12'd13,-12'd28,-12'd2,12'd61,12'd17,-12'd8,-12'd71,12'd1,-12'd41,-12'd7,-12'd34,12'd38,12'd61,-12'd22,12'd18,-12'd2,12'd5,-12'd5,12'd56,-12'd3,12'd43,12'd76,12'd5,-12'd28,12'd5,-12'd49,-12'd11,12'd24,-12'd3,-12'd5,12'd58,12'd2,12'd3,12'd18,-12'd45,12'd36,-12'd34,12'd15,-12'd29,-12'd32,-12'd35,-12'd32,12'd32,12'd27,12'd61,12'd9,12'd4,-12'd64,-12'd5,12'd52,12'd60,12'd29,12'd10,12'd58,-12'd37,12'd37,12'd47,12'd45,12'd35,-12'd22,12'd50,12'd6,12'd11,-12'd12,-12'd37,-12'd5,-12'd12,-12'd52,-12'd21,-12'd18,12'd35,-12'd6,-12'd60,12'd16,12'd13,-12'd31,-12'd20,-12'd47,-12'd16,-12'd11,-12'd15,-12'd38,12'd24,-12'd7,-12'd31,-12'd34,12'd44,-12'd12,12'd8,12'd21,-12'd33,12'd9,-12'd35,-12'd41,-12'd25,12'd28,12'd34,12'd24,12'd44,12'd25,-12'd11,-12'd7,-12'd28,-12'd1,12'd34,12'd29,-12'd21,-12'd18,-12'd13,-12'd20,12'd2,-12'd7,-12'd50,-12'd18,12'd43,12'd19,-12'd1,-12'd28,12'd12,-12'd42,-12'd15,12'd9,12'd25,-12'd51,-12'd39,-12'd21,12'd39,12'd37,-12'd15,-12'd27,-12'd4,-12'd42,-12'd45,-12'd30,-12'd17,-12'd18,12'd13,12'd14,12'd3,-12'd38,12'd36,12'd24,-12'd10,12'd32,-12'd11,12'd52,-12'd30,-12'd35,12'd39,-12'd34,12'd31,12'd55,-12'd31,-12'd19,-12'd3,-12'd8,-12'd32,-12'd66,12'd31,12'd11,12'd70,12'd20,-12'd28,-12'd5,12'd13,-12'd16,12'd11,-12'd25,-12'd2,12'd2,-12'd42,-12'd17,-12'd28,12'd3,-12'd24,12'd20,12'd29,-12'd45,12'd43,-12'd15,-12'd4,12'd63,12'd40,12'd30,-12'd7,-12'd35,-12'd1,12'd14,12'd26,-12'd51,-12'd29,12'd25,12'd0,12'd25,-12'd18,12'd16,-12'd22,-12'd35,12'd24,12'd14,12'd30,-12'd45,-12'd6,-12'd12,-12'd46,-12'd47,-12'd63,12'd7,-12'd37,12'd44,12'd29,-12'd24,12'd43,12'd12,-12'd5,-12'd17,12'd32,-12'd5,12'd15,12'd22,12'd16,-12'd18,-12'd17,-12'd29,-12'd1,12'd24,12'd59,-12'd62,-12'd6,12'd32,-12'd27,12'd72,-12'd19,-12'd1};

	clk = 0;
	#5 rst = 1;
	#10 rst = 0;
end

always
	#5 clk <= !clk;

endmodule

