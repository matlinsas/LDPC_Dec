`ifdef SIMULATION
    `include "cnu/cnu.v"
    `include "vnu/vnu.v"
    `include "check.v"
`endif

module ldpc_core(en, clk, rst, l/*, mtx*/, res, term, err);
parameter data_w = 6;
parameter mtx_w = 8;
parameter R = 24;
parameter C = 12;
parameter D = 96;
parameter N = 6;
localparam ext_w = log2(N);
localparam idx_w = 3;//log2(R);
localparam temp_w = data_w + ext_w;
localparam count_w = 5;

input clk, rst, en;
input [R*D*data_w-1:0] l;
//input [C*R*mtx_w-1:0] mtx;
output reg term;
output reg err;
output reg [R*D-1:0] res;

reg [count_w-1:0] count;

wire check;
wire [R*D-1:0] dec;

//check #(.mtx_w(mtx_w), .C(C), .R(R), .D(D)) CH (.dec(dec), .mtx(mtx), .res(check));
assign check = 1'b1;
always @(posedge clk) begin
	if(rst) begin
		res <= 0;
		err <= 0;
		count <= 0;
		term <= 1'b0;
    end else begin
        if(en) begin
            count <= count + 1'b1;
            if(count[count_w-1] || ~check) begin
                res <= dec;
				err <= check;
                term <= 1'b1;
            end
        end
    end
end

//------------------------------------------

function integer log2;
    input integer x;
    begin
        log2 = 0;
        while (x) begin
            log2 = log2 + 1;
            x = x>>1;
        end
    end
endfunction

//----------- Connections ----------------

wire [temp_w*6-1:0] c0ibus;
wire [data_w*6-1:0] c0obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU0 ( .en(en), .clk(clk), .rst(rst), .q(c0ibus), .r(c0obus));
wire [temp_w*6-1:0] c1ibus;
wire [data_w*6-1:0] c1obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1 ( .en(en), .clk(clk), .rst(rst), .q(c1ibus), .r(c1obus));
wire [temp_w*6-1:0] c2ibus;
wire [data_w*6-1:0] c2obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU2 ( .en(en), .clk(clk), .rst(rst), .q(c2ibus), .r(c2obus));
wire [temp_w*6-1:0] c3ibus;
wire [data_w*6-1:0] c3obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU3 ( .en(en), .clk(clk), .rst(rst), .q(c3ibus), .r(c3obus));
wire [temp_w*6-1:0] c4ibus;
wire [data_w*6-1:0] c4obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU4 ( .en(en), .clk(clk), .rst(rst), .q(c4ibus), .r(c4obus));
wire [temp_w*6-1:0] c5ibus;
wire [data_w*6-1:0] c5obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU5 ( .en(en), .clk(clk), .rst(rst), .q(c5ibus), .r(c5obus));
wire [temp_w*6-1:0] c6ibus;
wire [data_w*6-1:0] c6obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU6 ( .en(en), .clk(clk), .rst(rst), .q(c6ibus), .r(c6obus));
wire [temp_w*6-1:0] c7ibus;
wire [data_w*6-1:0] c7obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU7 ( .en(en), .clk(clk), .rst(rst), .q(c7ibus), .r(c7obus));
wire [temp_w*6-1:0] c8ibus;
wire [data_w*6-1:0] c8obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU8 ( .en(en), .clk(clk), .rst(rst), .q(c8ibus), .r(c8obus));
wire [temp_w*6-1:0] c9ibus;
wire [data_w*6-1:0] c9obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU9 ( .en(en), .clk(clk), .rst(rst), .q(c9ibus), .r(c9obus));
wire [temp_w*6-1:0] c10ibus;
wire [data_w*6-1:0] c10obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU10 ( .en(en), .clk(clk), .rst(rst), .q(c10ibus), .r(c10obus));
wire [temp_w*6-1:0] c11ibus;
wire [data_w*6-1:0] c11obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU11 ( .en(en), .clk(clk), .rst(rst), .q(c11ibus), .r(c11obus));
wire [temp_w*6-1:0] c12ibus;
wire [data_w*6-1:0] c12obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU12 ( .en(en), .clk(clk), .rst(rst), .q(c12ibus), .r(c12obus));
wire [temp_w*6-1:0] c13ibus;
wire [data_w*6-1:0] c13obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU13 ( .en(en), .clk(clk), .rst(rst), .q(c13ibus), .r(c13obus));
wire [temp_w*6-1:0] c14ibus;
wire [data_w*6-1:0] c14obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU14 ( .en(en), .clk(clk), .rst(rst), .q(c14ibus), .r(c14obus));
wire [temp_w*6-1:0] c15ibus;
wire [data_w*6-1:0] c15obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU15 ( .en(en), .clk(clk), .rst(rst), .q(c15ibus), .r(c15obus));
wire [temp_w*6-1:0] c16ibus;
wire [data_w*6-1:0] c16obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU16 ( .en(en), .clk(clk), .rst(rst), .q(c16ibus), .r(c16obus));
wire [temp_w*6-1:0] c17ibus;
wire [data_w*6-1:0] c17obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU17 ( .en(en), .clk(clk), .rst(rst), .q(c17ibus), .r(c17obus));
wire [temp_w*6-1:0] c18ibus;
wire [data_w*6-1:0] c18obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU18 ( .en(en), .clk(clk), .rst(rst), .q(c18ibus), .r(c18obus));
wire [temp_w*6-1:0] c19ibus;
wire [data_w*6-1:0] c19obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU19 ( .en(en), .clk(clk), .rst(rst), .q(c19ibus), .r(c19obus));
wire [temp_w*6-1:0] c20ibus;
wire [data_w*6-1:0] c20obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU20 ( .en(en), .clk(clk), .rst(rst), .q(c20ibus), .r(c20obus));
wire [temp_w*6-1:0] c21ibus;
wire [data_w*6-1:0] c21obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU21 ( .en(en), .clk(clk), .rst(rst), .q(c21ibus), .r(c21obus));
wire [temp_w*6-1:0] c22ibus;
wire [data_w*6-1:0] c22obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU22 ( .en(en), .clk(clk), .rst(rst), .q(c22ibus), .r(c22obus));
wire [temp_w*6-1:0] c23ibus;
wire [data_w*6-1:0] c23obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU23 ( .en(en), .clk(clk), .rst(rst), .q(c23ibus), .r(c23obus));
wire [temp_w*6-1:0] c24ibus;
wire [data_w*6-1:0] c24obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU24 ( .en(en), .clk(clk), .rst(rst), .q(c24ibus), .r(c24obus));
wire [temp_w*6-1:0] c25ibus;
wire [data_w*6-1:0] c25obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU25 ( .en(en), .clk(clk), .rst(rst), .q(c25ibus), .r(c25obus));
wire [temp_w*6-1:0] c26ibus;
wire [data_w*6-1:0] c26obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU26 ( .en(en), .clk(clk), .rst(rst), .q(c26ibus), .r(c26obus));
wire [temp_w*6-1:0] c27ibus;
wire [data_w*6-1:0] c27obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU27 ( .en(en), .clk(clk), .rst(rst), .q(c27ibus), .r(c27obus));
wire [temp_w*6-1:0] c28ibus;
wire [data_w*6-1:0] c28obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU28 ( .en(en), .clk(clk), .rst(rst), .q(c28ibus), .r(c28obus));
wire [temp_w*6-1:0] c29ibus;
wire [data_w*6-1:0] c29obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU29 ( .en(en), .clk(clk), .rst(rst), .q(c29ibus), .r(c29obus));
wire [temp_w*6-1:0] c30ibus;
wire [data_w*6-1:0] c30obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU30 ( .en(en), .clk(clk), .rst(rst), .q(c30ibus), .r(c30obus));
wire [temp_w*6-1:0] c31ibus;
wire [data_w*6-1:0] c31obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU31 ( .en(en), .clk(clk), .rst(rst), .q(c31ibus), .r(c31obus));
wire [temp_w*6-1:0] c32ibus;
wire [data_w*6-1:0] c32obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU32 ( .en(en), .clk(clk), .rst(rst), .q(c32ibus), .r(c32obus));
wire [temp_w*6-1:0] c33ibus;
wire [data_w*6-1:0] c33obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU33 ( .en(en), .clk(clk), .rst(rst), .q(c33ibus), .r(c33obus));
wire [temp_w*6-1:0] c34ibus;
wire [data_w*6-1:0] c34obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU34 ( .en(en), .clk(clk), .rst(rst), .q(c34ibus), .r(c34obus));
wire [temp_w*6-1:0] c35ibus;
wire [data_w*6-1:0] c35obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU35 ( .en(en), .clk(clk), .rst(rst), .q(c35ibus), .r(c35obus));
wire [temp_w*6-1:0] c36ibus;
wire [data_w*6-1:0] c36obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU36 ( .en(en), .clk(clk), .rst(rst), .q(c36ibus), .r(c36obus));
wire [temp_w*6-1:0] c37ibus;
wire [data_w*6-1:0] c37obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU37 ( .en(en), .clk(clk), .rst(rst), .q(c37ibus), .r(c37obus));
wire [temp_w*6-1:0] c38ibus;
wire [data_w*6-1:0] c38obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU38 ( .en(en), .clk(clk), .rst(rst), .q(c38ibus), .r(c38obus));
wire [temp_w*6-1:0] c39ibus;
wire [data_w*6-1:0] c39obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU39 ( .en(en), .clk(clk), .rst(rst), .q(c39ibus), .r(c39obus));
wire [temp_w*6-1:0] c40ibus;
wire [data_w*6-1:0] c40obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU40 ( .en(en), .clk(clk), .rst(rst), .q(c40ibus), .r(c40obus));
wire [temp_w*6-1:0] c41ibus;
wire [data_w*6-1:0] c41obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU41 ( .en(en), .clk(clk), .rst(rst), .q(c41ibus), .r(c41obus));
wire [temp_w*6-1:0] c42ibus;
wire [data_w*6-1:0] c42obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU42 ( .en(en), .clk(clk), .rst(rst), .q(c42ibus), .r(c42obus));
wire [temp_w*6-1:0] c43ibus;
wire [data_w*6-1:0] c43obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU43 ( .en(en), .clk(clk), .rst(rst), .q(c43ibus), .r(c43obus));
wire [temp_w*6-1:0] c44ibus;
wire [data_w*6-1:0] c44obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU44 ( .en(en), .clk(clk), .rst(rst), .q(c44ibus), .r(c44obus));
wire [temp_w*6-1:0] c45ibus;
wire [data_w*6-1:0] c45obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU45 ( .en(en), .clk(clk), .rst(rst), .q(c45ibus), .r(c45obus));
wire [temp_w*6-1:0] c46ibus;
wire [data_w*6-1:0] c46obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU46 ( .en(en), .clk(clk), .rst(rst), .q(c46ibus), .r(c46obus));
wire [temp_w*6-1:0] c47ibus;
wire [data_w*6-1:0] c47obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU47 ( .en(en), .clk(clk), .rst(rst), .q(c47ibus), .r(c47obus));
wire [temp_w*6-1:0] c48ibus;
wire [data_w*6-1:0] c48obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU48 ( .en(en), .clk(clk), .rst(rst), .q(c48ibus), .r(c48obus));
wire [temp_w*6-1:0] c49ibus;
wire [data_w*6-1:0] c49obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU49 ( .en(en), .clk(clk), .rst(rst), .q(c49ibus), .r(c49obus));
wire [temp_w*6-1:0] c50ibus;
wire [data_w*6-1:0] c50obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU50 ( .en(en), .clk(clk), .rst(rst), .q(c50ibus), .r(c50obus));
wire [temp_w*6-1:0] c51ibus;
wire [data_w*6-1:0] c51obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU51 ( .en(en), .clk(clk), .rst(rst), .q(c51ibus), .r(c51obus));
wire [temp_w*6-1:0] c52ibus;
wire [data_w*6-1:0] c52obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU52 ( .en(en), .clk(clk), .rst(rst), .q(c52ibus), .r(c52obus));
wire [temp_w*6-1:0] c53ibus;
wire [data_w*6-1:0] c53obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU53 ( .en(en), .clk(clk), .rst(rst), .q(c53ibus), .r(c53obus));
wire [temp_w*6-1:0] c54ibus;
wire [data_w*6-1:0] c54obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU54 ( .en(en), .clk(clk), .rst(rst), .q(c54ibus), .r(c54obus));
wire [temp_w*6-1:0] c55ibus;
wire [data_w*6-1:0] c55obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU55 ( .en(en), .clk(clk), .rst(rst), .q(c55ibus), .r(c55obus));
wire [temp_w*6-1:0] c56ibus;
wire [data_w*6-1:0] c56obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU56 ( .en(en), .clk(clk), .rst(rst), .q(c56ibus), .r(c56obus));
wire [temp_w*6-1:0] c57ibus;
wire [data_w*6-1:0] c57obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU57 ( .en(en), .clk(clk), .rst(rst), .q(c57ibus), .r(c57obus));
wire [temp_w*6-1:0] c58ibus;
wire [data_w*6-1:0] c58obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU58 ( .en(en), .clk(clk), .rst(rst), .q(c58ibus), .r(c58obus));
wire [temp_w*6-1:0] c59ibus;
wire [data_w*6-1:0] c59obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU59 ( .en(en), .clk(clk), .rst(rst), .q(c59ibus), .r(c59obus));
wire [temp_w*6-1:0] c60ibus;
wire [data_w*6-1:0] c60obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU60 ( .en(en), .clk(clk), .rst(rst), .q(c60ibus), .r(c60obus));
wire [temp_w*6-1:0] c61ibus;
wire [data_w*6-1:0] c61obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU61 ( .en(en), .clk(clk), .rst(rst), .q(c61ibus), .r(c61obus));
wire [temp_w*6-1:0] c62ibus;
wire [data_w*6-1:0] c62obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU62 ( .en(en), .clk(clk), .rst(rst), .q(c62ibus), .r(c62obus));
wire [temp_w*6-1:0] c63ibus;
wire [data_w*6-1:0] c63obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU63 ( .en(en), .clk(clk), .rst(rst), .q(c63ibus), .r(c63obus));
wire [temp_w*6-1:0] c64ibus;
wire [data_w*6-1:0] c64obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU64 ( .en(en), .clk(clk), .rst(rst), .q(c64ibus), .r(c64obus));
wire [temp_w*6-1:0] c65ibus;
wire [data_w*6-1:0] c65obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU65 ( .en(en), .clk(clk), .rst(rst), .q(c65ibus), .r(c65obus));
wire [temp_w*6-1:0] c66ibus;
wire [data_w*6-1:0] c66obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU66 ( .en(en), .clk(clk), .rst(rst), .q(c66ibus), .r(c66obus));
wire [temp_w*6-1:0] c67ibus;
wire [data_w*6-1:0] c67obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU67 ( .en(en), .clk(clk), .rst(rst), .q(c67ibus), .r(c67obus));
wire [temp_w*6-1:0] c68ibus;
wire [data_w*6-1:0] c68obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU68 ( .en(en), .clk(clk), .rst(rst), .q(c68ibus), .r(c68obus));
wire [temp_w*6-1:0] c69ibus;
wire [data_w*6-1:0] c69obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU69 ( .en(en), .clk(clk), .rst(rst), .q(c69ibus), .r(c69obus));
wire [temp_w*6-1:0] c70ibus;
wire [data_w*6-1:0] c70obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU70 ( .en(en), .clk(clk), .rst(rst), .q(c70ibus), .r(c70obus));
wire [temp_w*6-1:0] c71ibus;
wire [data_w*6-1:0] c71obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU71 ( .en(en), .clk(clk), .rst(rst), .q(c71ibus), .r(c71obus));
wire [temp_w*6-1:0] c72ibus;
wire [data_w*6-1:0] c72obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU72 ( .en(en), .clk(clk), .rst(rst), .q(c72ibus), .r(c72obus));
wire [temp_w*6-1:0] c73ibus;
wire [data_w*6-1:0] c73obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU73 ( .en(en), .clk(clk), .rst(rst), .q(c73ibus), .r(c73obus));
wire [temp_w*6-1:0] c74ibus;
wire [data_w*6-1:0] c74obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU74 ( .en(en), .clk(clk), .rst(rst), .q(c74ibus), .r(c74obus));
wire [temp_w*6-1:0] c75ibus;
wire [data_w*6-1:0] c75obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU75 ( .en(en), .clk(clk), .rst(rst), .q(c75ibus), .r(c75obus));
wire [temp_w*6-1:0] c76ibus;
wire [data_w*6-1:0] c76obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU76 ( .en(en), .clk(clk), .rst(rst), .q(c76ibus), .r(c76obus));
wire [temp_w*6-1:0] c77ibus;
wire [data_w*6-1:0] c77obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU77 ( .en(en), .clk(clk), .rst(rst), .q(c77ibus), .r(c77obus));
wire [temp_w*6-1:0] c78ibus;
wire [data_w*6-1:0] c78obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU78 ( .en(en), .clk(clk), .rst(rst), .q(c78ibus), .r(c78obus));
wire [temp_w*6-1:0] c79ibus;
wire [data_w*6-1:0] c79obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU79 ( .en(en), .clk(clk), .rst(rst), .q(c79ibus), .r(c79obus));
wire [temp_w*6-1:0] c80ibus;
wire [data_w*6-1:0] c80obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU80 ( .en(en), .clk(clk), .rst(rst), .q(c80ibus), .r(c80obus));
wire [temp_w*6-1:0] c81ibus;
wire [data_w*6-1:0] c81obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU81 ( .en(en), .clk(clk), .rst(rst), .q(c81ibus), .r(c81obus));
wire [temp_w*6-1:0] c82ibus;
wire [data_w*6-1:0] c82obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU82 ( .en(en), .clk(clk), .rst(rst), .q(c82ibus), .r(c82obus));
wire [temp_w*6-1:0] c83ibus;
wire [data_w*6-1:0] c83obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU83 ( .en(en), .clk(clk), .rst(rst), .q(c83ibus), .r(c83obus));
wire [temp_w*6-1:0] c84ibus;
wire [data_w*6-1:0] c84obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU84 ( .en(en), .clk(clk), .rst(rst), .q(c84ibus), .r(c84obus));
wire [temp_w*6-1:0] c85ibus;
wire [data_w*6-1:0] c85obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU85 ( .en(en), .clk(clk), .rst(rst), .q(c85ibus), .r(c85obus));
wire [temp_w*6-1:0] c86ibus;
wire [data_w*6-1:0] c86obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU86 ( .en(en), .clk(clk), .rst(rst), .q(c86ibus), .r(c86obus));
wire [temp_w*6-1:0] c87ibus;
wire [data_w*6-1:0] c87obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU87 ( .en(en), .clk(clk), .rst(rst), .q(c87ibus), .r(c87obus));
wire [temp_w*6-1:0] c88ibus;
wire [data_w*6-1:0] c88obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU88 ( .en(en), .clk(clk), .rst(rst), .q(c88ibus), .r(c88obus));
wire [temp_w*6-1:0] c89ibus;
wire [data_w*6-1:0] c89obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU89 ( .en(en), .clk(clk), .rst(rst), .q(c89ibus), .r(c89obus));
wire [temp_w*6-1:0] c90ibus;
wire [data_w*6-1:0] c90obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU90 ( .en(en), .clk(clk), .rst(rst), .q(c90ibus), .r(c90obus));
wire [temp_w*6-1:0] c91ibus;
wire [data_w*6-1:0] c91obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU91 ( .en(en), .clk(clk), .rst(rst), .q(c91ibus), .r(c91obus));
wire [temp_w*6-1:0] c92ibus;
wire [data_w*6-1:0] c92obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU92 ( .en(en), .clk(clk), .rst(rst), .q(c92ibus), .r(c92obus));
wire [temp_w*6-1:0] c93ibus;
wire [data_w*6-1:0] c93obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU93 ( .en(en), .clk(clk), .rst(rst), .q(c93ibus), .r(c93obus));
wire [temp_w*6-1:0] c94ibus;
wire [data_w*6-1:0] c94obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU94 ( .en(en), .clk(clk), .rst(rst), .q(c94ibus), .r(c94obus));
wire [temp_w*6-1:0] c95ibus;
wire [data_w*6-1:0] c95obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU95 ( .en(en), .clk(clk), .rst(rst), .q(c95ibus), .r(c95obus));
wire [temp_w*7-1:0] c96ibus;
wire [data_w*7-1:0] c96obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU96 ( .en(en), .clk(clk), .rst(rst), .q(c96ibus), .r(c96obus));
wire [temp_w*7-1:0] c97ibus;
wire [data_w*7-1:0] c97obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU97 ( .en(en), .clk(clk), .rst(rst), .q(c97ibus), .r(c97obus));
wire [temp_w*7-1:0] c98ibus;
wire [data_w*7-1:0] c98obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU98 ( .en(en), .clk(clk), .rst(rst), .q(c98ibus), .r(c98obus));
wire [temp_w*7-1:0] c99ibus;
wire [data_w*7-1:0] c99obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU99 ( .en(en), .clk(clk), .rst(rst), .q(c99ibus), .r(c99obus));
wire [temp_w*7-1:0] c100ibus;
wire [data_w*7-1:0] c100obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU100 ( .en(en), .clk(clk), .rst(rst), .q(c100ibus), .r(c100obus));
wire [temp_w*7-1:0] c101ibus;
wire [data_w*7-1:0] c101obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU101 ( .en(en), .clk(clk), .rst(rst), .q(c101ibus), .r(c101obus));
wire [temp_w*7-1:0] c102ibus;
wire [data_w*7-1:0] c102obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU102 ( .en(en), .clk(clk), .rst(rst), .q(c102ibus), .r(c102obus));
wire [temp_w*7-1:0] c103ibus;
wire [data_w*7-1:0] c103obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU103 ( .en(en), .clk(clk), .rst(rst), .q(c103ibus), .r(c103obus));
wire [temp_w*7-1:0] c104ibus;
wire [data_w*7-1:0] c104obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU104 ( .en(en), .clk(clk), .rst(rst), .q(c104ibus), .r(c104obus));
wire [temp_w*7-1:0] c105ibus;
wire [data_w*7-1:0] c105obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU105 ( .en(en), .clk(clk), .rst(rst), .q(c105ibus), .r(c105obus));
wire [temp_w*7-1:0] c106ibus;
wire [data_w*7-1:0] c106obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU106 ( .en(en), .clk(clk), .rst(rst), .q(c106ibus), .r(c106obus));
wire [temp_w*7-1:0] c107ibus;
wire [data_w*7-1:0] c107obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU107 ( .en(en), .clk(clk), .rst(rst), .q(c107ibus), .r(c107obus));
wire [temp_w*7-1:0] c108ibus;
wire [data_w*7-1:0] c108obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU108 ( .en(en), .clk(clk), .rst(rst), .q(c108ibus), .r(c108obus));
wire [temp_w*7-1:0] c109ibus;
wire [data_w*7-1:0] c109obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU109 ( .en(en), .clk(clk), .rst(rst), .q(c109ibus), .r(c109obus));
wire [temp_w*7-1:0] c110ibus;
wire [data_w*7-1:0] c110obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU110 ( .en(en), .clk(clk), .rst(rst), .q(c110ibus), .r(c110obus));
wire [temp_w*7-1:0] c111ibus;
wire [data_w*7-1:0] c111obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU111 ( .en(en), .clk(clk), .rst(rst), .q(c111ibus), .r(c111obus));
wire [temp_w*7-1:0] c112ibus;
wire [data_w*7-1:0] c112obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU112 ( .en(en), .clk(clk), .rst(rst), .q(c112ibus), .r(c112obus));
wire [temp_w*7-1:0] c113ibus;
wire [data_w*7-1:0] c113obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU113 ( .en(en), .clk(clk), .rst(rst), .q(c113ibus), .r(c113obus));
wire [temp_w*7-1:0] c114ibus;
wire [data_w*7-1:0] c114obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU114 ( .en(en), .clk(clk), .rst(rst), .q(c114ibus), .r(c114obus));
wire [temp_w*7-1:0] c115ibus;
wire [data_w*7-1:0] c115obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU115 ( .en(en), .clk(clk), .rst(rst), .q(c115ibus), .r(c115obus));
wire [temp_w*7-1:0] c116ibus;
wire [data_w*7-1:0] c116obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU116 ( .en(en), .clk(clk), .rst(rst), .q(c116ibus), .r(c116obus));
wire [temp_w*7-1:0] c117ibus;
wire [data_w*7-1:0] c117obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU117 ( .en(en), .clk(clk), .rst(rst), .q(c117ibus), .r(c117obus));
wire [temp_w*7-1:0] c118ibus;
wire [data_w*7-1:0] c118obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU118 ( .en(en), .clk(clk), .rst(rst), .q(c118ibus), .r(c118obus));
wire [temp_w*7-1:0] c119ibus;
wire [data_w*7-1:0] c119obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU119 ( .en(en), .clk(clk), .rst(rst), .q(c119ibus), .r(c119obus));
wire [temp_w*7-1:0] c120ibus;
wire [data_w*7-1:0] c120obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU120 ( .en(en), .clk(clk), .rst(rst), .q(c120ibus), .r(c120obus));
wire [temp_w*7-1:0] c121ibus;
wire [data_w*7-1:0] c121obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU121 ( .en(en), .clk(clk), .rst(rst), .q(c121ibus), .r(c121obus));
wire [temp_w*7-1:0] c122ibus;
wire [data_w*7-1:0] c122obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU122 ( .en(en), .clk(clk), .rst(rst), .q(c122ibus), .r(c122obus));
wire [temp_w*7-1:0] c123ibus;
wire [data_w*7-1:0] c123obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU123 ( .en(en), .clk(clk), .rst(rst), .q(c123ibus), .r(c123obus));
wire [temp_w*7-1:0] c124ibus;
wire [data_w*7-1:0] c124obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU124 ( .en(en), .clk(clk), .rst(rst), .q(c124ibus), .r(c124obus));
wire [temp_w*7-1:0] c125ibus;
wire [data_w*7-1:0] c125obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU125 ( .en(en), .clk(clk), .rst(rst), .q(c125ibus), .r(c125obus));
wire [temp_w*7-1:0] c126ibus;
wire [data_w*7-1:0] c126obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU126 ( .en(en), .clk(clk), .rst(rst), .q(c126ibus), .r(c126obus));
wire [temp_w*7-1:0] c127ibus;
wire [data_w*7-1:0] c127obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU127 ( .en(en), .clk(clk), .rst(rst), .q(c127ibus), .r(c127obus));
wire [temp_w*7-1:0] c128ibus;
wire [data_w*7-1:0] c128obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU128 ( .en(en), .clk(clk), .rst(rst), .q(c128ibus), .r(c128obus));
wire [temp_w*7-1:0] c129ibus;
wire [data_w*7-1:0] c129obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU129 ( .en(en), .clk(clk), .rst(rst), .q(c129ibus), .r(c129obus));
wire [temp_w*7-1:0] c130ibus;
wire [data_w*7-1:0] c130obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU130 ( .en(en), .clk(clk), .rst(rst), .q(c130ibus), .r(c130obus));
wire [temp_w*7-1:0] c131ibus;
wire [data_w*7-1:0] c131obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU131 ( .en(en), .clk(clk), .rst(rst), .q(c131ibus), .r(c131obus));
wire [temp_w*7-1:0] c132ibus;
wire [data_w*7-1:0] c132obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU132 ( .en(en), .clk(clk), .rst(rst), .q(c132ibus), .r(c132obus));
wire [temp_w*7-1:0] c133ibus;
wire [data_w*7-1:0] c133obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU133 ( .en(en), .clk(clk), .rst(rst), .q(c133ibus), .r(c133obus));
wire [temp_w*7-1:0] c134ibus;
wire [data_w*7-1:0] c134obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU134 ( .en(en), .clk(clk), .rst(rst), .q(c134ibus), .r(c134obus));
wire [temp_w*7-1:0] c135ibus;
wire [data_w*7-1:0] c135obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU135 ( .en(en), .clk(clk), .rst(rst), .q(c135ibus), .r(c135obus));
wire [temp_w*7-1:0] c136ibus;
wire [data_w*7-1:0] c136obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU136 ( .en(en), .clk(clk), .rst(rst), .q(c136ibus), .r(c136obus));
wire [temp_w*7-1:0] c137ibus;
wire [data_w*7-1:0] c137obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU137 ( .en(en), .clk(clk), .rst(rst), .q(c137ibus), .r(c137obus));
wire [temp_w*7-1:0] c138ibus;
wire [data_w*7-1:0] c138obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU138 ( .en(en), .clk(clk), .rst(rst), .q(c138ibus), .r(c138obus));
wire [temp_w*7-1:0] c139ibus;
wire [data_w*7-1:0] c139obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU139 ( .en(en), .clk(clk), .rst(rst), .q(c139ibus), .r(c139obus));
wire [temp_w*7-1:0] c140ibus;
wire [data_w*7-1:0] c140obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU140 ( .en(en), .clk(clk), .rst(rst), .q(c140ibus), .r(c140obus));
wire [temp_w*7-1:0] c141ibus;
wire [data_w*7-1:0] c141obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU141 ( .en(en), .clk(clk), .rst(rst), .q(c141ibus), .r(c141obus));
wire [temp_w*7-1:0] c142ibus;
wire [data_w*7-1:0] c142obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU142 ( .en(en), .clk(clk), .rst(rst), .q(c142ibus), .r(c142obus));
wire [temp_w*7-1:0] c143ibus;
wire [data_w*7-1:0] c143obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU143 ( .en(en), .clk(clk), .rst(rst), .q(c143ibus), .r(c143obus));
wire [temp_w*7-1:0] c144ibus;
wire [data_w*7-1:0] c144obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU144 ( .en(en), .clk(clk), .rst(rst), .q(c144ibus), .r(c144obus));
wire [temp_w*7-1:0] c145ibus;
wire [data_w*7-1:0] c145obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU145 ( .en(en), .clk(clk), .rst(rst), .q(c145ibus), .r(c145obus));
wire [temp_w*7-1:0] c146ibus;
wire [data_w*7-1:0] c146obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU146 ( .en(en), .clk(clk), .rst(rst), .q(c146ibus), .r(c146obus));
wire [temp_w*7-1:0] c147ibus;
wire [data_w*7-1:0] c147obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU147 ( .en(en), .clk(clk), .rst(rst), .q(c147ibus), .r(c147obus));
wire [temp_w*7-1:0] c148ibus;
wire [data_w*7-1:0] c148obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU148 ( .en(en), .clk(clk), .rst(rst), .q(c148ibus), .r(c148obus));
wire [temp_w*7-1:0] c149ibus;
wire [data_w*7-1:0] c149obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU149 ( .en(en), .clk(clk), .rst(rst), .q(c149ibus), .r(c149obus));
wire [temp_w*7-1:0] c150ibus;
wire [data_w*7-1:0] c150obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU150 ( .en(en), .clk(clk), .rst(rst), .q(c150ibus), .r(c150obus));
wire [temp_w*7-1:0] c151ibus;
wire [data_w*7-1:0] c151obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU151 ( .en(en), .clk(clk), .rst(rst), .q(c151ibus), .r(c151obus));
wire [temp_w*7-1:0] c152ibus;
wire [data_w*7-1:0] c152obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU152 ( .en(en), .clk(clk), .rst(rst), .q(c152ibus), .r(c152obus));
wire [temp_w*7-1:0] c153ibus;
wire [data_w*7-1:0] c153obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU153 ( .en(en), .clk(clk), .rst(rst), .q(c153ibus), .r(c153obus));
wire [temp_w*7-1:0] c154ibus;
wire [data_w*7-1:0] c154obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU154 ( .en(en), .clk(clk), .rst(rst), .q(c154ibus), .r(c154obus));
wire [temp_w*7-1:0] c155ibus;
wire [data_w*7-1:0] c155obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU155 ( .en(en), .clk(clk), .rst(rst), .q(c155ibus), .r(c155obus));
wire [temp_w*7-1:0] c156ibus;
wire [data_w*7-1:0] c156obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU156 ( .en(en), .clk(clk), .rst(rst), .q(c156ibus), .r(c156obus));
wire [temp_w*7-1:0] c157ibus;
wire [data_w*7-1:0] c157obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU157 ( .en(en), .clk(clk), .rst(rst), .q(c157ibus), .r(c157obus));
wire [temp_w*7-1:0] c158ibus;
wire [data_w*7-1:0] c158obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU158 ( .en(en), .clk(clk), .rst(rst), .q(c158ibus), .r(c158obus));
wire [temp_w*7-1:0] c159ibus;
wire [data_w*7-1:0] c159obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU159 ( .en(en), .clk(clk), .rst(rst), .q(c159ibus), .r(c159obus));
wire [temp_w*7-1:0] c160ibus;
wire [data_w*7-1:0] c160obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU160 ( .en(en), .clk(clk), .rst(rst), .q(c160ibus), .r(c160obus));
wire [temp_w*7-1:0] c161ibus;
wire [data_w*7-1:0] c161obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU161 ( .en(en), .clk(clk), .rst(rst), .q(c161ibus), .r(c161obus));
wire [temp_w*7-1:0] c162ibus;
wire [data_w*7-1:0] c162obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU162 ( .en(en), .clk(clk), .rst(rst), .q(c162ibus), .r(c162obus));
wire [temp_w*7-1:0] c163ibus;
wire [data_w*7-1:0] c163obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU163 ( .en(en), .clk(clk), .rst(rst), .q(c163ibus), .r(c163obus));
wire [temp_w*7-1:0] c164ibus;
wire [data_w*7-1:0] c164obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU164 ( .en(en), .clk(clk), .rst(rst), .q(c164ibus), .r(c164obus));
wire [temp_w*7-1:0] c165ibus;
wire [data_w*7-1:0] c165obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU165 ( .en(en), .clk(clk), .rst(rst), .q(c165ibus), .r(c165obus));
wire [temp_w*7-1:0] c166ibus;
wire [data_w*7-1:0] c166obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU166 ( .en(en), .clk(clk), .rst(rst), .q(c166ibus), .r(c166obus));
wire [temp_w*7-1:0] c167ibus;
wire [data_w*7-1:0] c167obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU167 ( .en(en), .clk(clk), .rst(rst), .q(c167ibus), .r(c167obus));
wire [temp_w*7-1:0] c168ibus;
wire [data_w*7-1:0] c168obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU168 ( .en(en), .clk(clk), .rst(rst), .q(c168ibus), .r(c168obus));
wire [temp_w*7-1:0] c169ibus;
wire [data_w*7-1:0] c169obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU169 ( .en(en), .clk(clk), .rst(rst), .q(c169ibus), .r(c169obus));
wire [temp_w*7-1:0] c170ibus;
wire [data_w*7-1:0] c170obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU170 ( .en(en), .clk(clk), .rst(rst), .q(c170ibus), .r(c170obus));
wire [temp_w*7-1:0] c171ibus;
wire [data_w*7-1:0] c171obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU171 ( .en(en), .clk(clk), .rst(rst), .q(c171ibus), .r(c171obus));
wire [temp_w*7-1:0] c172ibus;
wire [data_w*7-1:0] c172obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU172 ( .en(en), .clk(clk), .rst(rst), .q(c172ibus), .r(c172obus));
wire [temp_w*7-1:0] c173ibus;
wire [data_w*7-1:0] c173obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU173 ( .en(en), .clk(clk), .rst(rst), .q(c173ibus), .r(c173obus));
wire [temp_w*7-1:0] c174ibus;
wire [data_w*7-1:0] c174obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU174 ( .en(en), .clk(clk), .rst(rst), .q(c174ibus), .r(c174obus));
wire [temp_w*7-1:0] c175ibus;
wire [data_w*7-1:0] c175obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU175 ( .en(en), .clk(clk), .rst(rst), .q(c175ibus), .r(c175obus));
wire [temp_w*7-1:0] c176ibus;
wire [data_w*7-1:0] c176obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU176 ( .en(en), .clk(clk), .rst(rst), .q(c176ibus), .r(c176obus));
wire [temp_w*7-1:0] c177ibus;
wire [data_w*7-1:0] c177obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU177 ( .en(en), .clk(clk), .rst(rst), .q(c177ibus), .r(c177obus));
wire [temp_w*7-1:0] c178ibus;
wire [data_w*7-1:0] c178obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU178 ( .en(en), .clk(clk), .rst(rst), .q(c178ibus), .r(c178obus));
wire [temp_w*7-1:0] c179ibus;
wire [data_w*7-1:0] c179obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU179 ( .en(en), .clk(clk), .rst(rst), .q(c179ibus), .r(c179obus));
wire [temp_w*7-1:0] c180ibus;
wire [data_w*7-1:0] c180obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU180 ( .en(en), .clk(clk), .rst(rst), .q(c180ibus), .r(c180obus));
wire [temp_w*7-1:0] c181ibus;
wire [data_w*7-1:0] c181obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU181 ( .en(en), .clk(clk), .rst(rst), .q(c181ibus), .r(c181obus));
wire [temp_w*7-1:0] c182ibus;
wire [data_w*7-1:0] c182obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU182 ( .en(en), .clk(clk), .rst(rst), .q(c182ibus), .r(c182obus));
wire [temp_w*7-1:0] c183ibus;
wire [data_w*7-1:0] c183obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU183 ( .en(en), .clk(clk), .rst(rst), .q(c183ibus), .r(c183obus));
wire [temp_w*7-1:0] c184ibus;
wire [data_w*7-1:0] c184obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU184 ( .en(en), .clk(clk), .rst(rst), .q(c184ibus), .r(c184obus));
wire [temp_w*7-1:0] c185ibus;
wire [data_w*7-1:0] c185obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU185 ( .en(en), .clk(clk), .rst(rst), .q(c185ibus), .r(c185obus));
wire [temp_w*7-1:0] c186ibus;
wire [data_w*7-1:0] c186obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU186 ( .en(en), .clk(clk), .rst(rst), .q(c186ibus), .r(c186obus));
wire [temp_w*7-1:0] c187ibus;
wire [data_w*7-1:0] c187obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU187 ( .en(en), .clk(clk), .rst(rst), .q(c187ibus), .r(c187obus));
wire [temp_w*7-1:0] c188ibus;
wire [data_w*7-1:0] c188obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU188 ( .en(en), .clk(clk), .rst(rst), .q(c188ibus), .r(c188obus));
wire [temp_w*7-1:0] c189ibus;
wire [data_w*7-1:0] c189obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU189 ( .en(en), .clk(clk), .rst(rst), .q(c189ibus), .r(c189obus));
wire [temp_w*7-1:0] c190ibus;
wire [data_w*7-1:0] c190obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU190 ( .en(en), .clk(clk), .rst(rst), .q(c190ibus), .r(c190obus));
wire [temp_w*7-1:0] c191ibus;
wire [data_w*7-1:0] c191obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU191 ( .en(en), .clk(clk), .rst(rst), .q(c191ibus), .r(c191obus));
wire [temp_w*7-1:0] c192ibus;
wire [data_w*7-1:0] c192obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU192 ( .en(en), .clk(clk), .rst(rst), .q(c192ibus), .r(c192obus));
wire [temp_w*7-1:0] c193ibus;
wire [data_w*7-1:0] c193obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU193 ( .en(en), .clk(clk), .rst(rst), .q(c193ibus), .r(c193obus));
wire [temp_w*7-1:0] c194ibus;
wire [data_w*7-1:0] c194obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU194 ( .en(en), .clk(clk), .rst(rst), .q(c194ibus), .r(c194obus));
wire [temp_w*7-1:0] c195ibus;
wire [data_w*7-1:0] c195obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU195 ( .en(en), .clk(clk), .rst(rst), .q(c195ibus), .r(c195obus));
wire [temp_w*7-1:0] c196ibus;
wire [data_w*7-1:0] c196obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU196 ( .en(en), .clk(clk), .rst(rst), .q(c196ibus), .r(c196obus));
wire [temp_w*7-1:0] c197ibus;
wire [data_w*7-1:0] c197obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU197 ( .en(en), .clk(clk), .rst(rst), .q(c197ibus), .r(c197obus));
wire [temp_w*7-1:0] c198ibus;
wire [data_w*7-1:0] c198obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU198 ( .en(en), .clk(clk), .rst(rst), .q(c198ibus), .r(c198obus));
wire [temp_w*7-1:0] c199ibus;
wire [data_w*7-1:0] c199obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU199 ( .en(en), .clk(clk), .rst(rst), .q(c199ibus), .r(c199obus));
wire [temp_w*7-1:0] c200ibus;
wire [data_w*7-1:0] c200obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU200 ( .en(en), .clk(clk), .rst(rst), .q(c200ibus), .r(c200obus));
wire [temp_w*7-1:0] c201ibus;
wire [data_w*7-1:0] c201obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU201 ( .en(en), .clk(clk), .rst(rst), .q(c201ibus), .r(c201obus));
wire [temp_w*7-1:0] c202ibus;
wire [data_w*7-1:0] c202obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU202 ( .en(en), .clk(clk), .rst(rst), .q(c202ibus), .r(c202obus));
wire [temp_w*7-1:0] c203ibus;
wire [data_w*7-1:0] c203obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU203 ( .en(en), .clk(clk), .rst(rst), .q(c203ibus), .r(c203obus));
wire [temp_w*7-1:0] c204ibus;
wire [data_w*7-1:0] c204obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU204 ( .en(en), .clk(clk), .rst(rst), .q(c204ibus), .r(c204obus));
wire [temp_w*7-1:0] c205ibus;
wire [data_w*7-1:0] c205obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU205 ( .en(en), .clk(clk), .rst(rst), .q(c205ibus), .r(c205obus));
wire [temp_w*7-1:0] c206ibus;
wire [data_w*7-1:0] c206obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU206 ( .en(en), .clk(clk), .rst(rst), .q(c206ibus), .r(c206obus));
wire [temp_w*7-1:0] c207ibus;
wire [data_w*7-1:0] c207obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU207 ( .en(en), .clk(clk), .rst(rst), .q(c207ibus), .r(c207obus));
wire [temp_w*7-1:0] c208ibus;
wire [data_w*7-1:0] c208obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU208 ( .en(en), .clk(clk), .rst(rst), .q(c208ibus), .r(c208obus));
wire [temp_w*7-1:0] c209ibus;
wire [data_w*7-1:0] c209obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU209 ( .en(en), .clk(clk), .rst(rst), .q(c209ibus), .r(c209obus));
wire [temp_w*7-1:0] c210ibus;
wire [data_w*7-1:0] c210obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU210 ( .en(en), .clk(clk), .rst(rst), .q(c210ibus), .r(c210obus));
wire [temp_w*7-1:0] c211ibus;
wire [data_w*7-1:0] c211obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU211 ( .en(en), .clk(clk), .rst(rst), .q(c211ibus), .r(c211obus));
wire [temp_w*7-1:0] c212ibus;
wire [data_w*7-1:0] c212obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU212 ( .en(en), .clk(clk), .rst(rst), .q(c212ibus), .r(c212obus));
wire [temp_w*7-1:0] c213ibus;
wire [data_w*7-1:0] c213obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU213 ( .en(en), .clk(clk), .rst(rst), .q(c213ibus), .r(c213obus));
wire [temp_w*7-1:0] c214ibus;
wire [data_w*7-1:0] c214obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU214 ( .en(en), .clk(clk), .rst(rst), .q(c214ibus), .r(c214obus));
wire [temp_w*7-1:0] c215ibus;
wire [data_w*7-1:0] c215obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU215 ( .en(en), .clk(clk), .rst(rst), .q(c215ibus), .r(c215obus));
wire [temp_w*7-1:0] c216ibus;
wire [data_w*7-1:0] c216obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU216 ( .en(en), .clk(clk), .rst(rst), .q(c216ibus), .r(c216obus));
wire [temp_w*7-1:0] c217ibus;
wire [data_w*7-1:0] c217obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU217 ( .en(en), .clk(clk), .rst(rst), .q(c217ibus), .r(c217obus));
wire [temp_w*7-1:0] c218ibus;
wire [data_w*7-1:0] c218obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU218 ( .en(en), .clk(clk), .rst(rst), .q(c218ibus), .r(c218obus));
wire [temp_w*7-1:0] c219ibus;
wire [data_w*7-1:0] c219obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU219 ( .en(en), .clk(clk), .rst(rst), .q(c219ibus), .r(c219obus));
wire [temp_w*7-1:0] c220ibus;
wire [data_w*7-1:0] c220obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU220 ( .en(en), .clk(clk), .rst(rst), .q(c220ibus), .r(c220obus));
wire [temp_w*7-1:0] c221ibus;
wire [data_w*7-1:0] c221obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU221 ( .en(en), .clk(clk), .rst(rst), .q(c221ibus), .r(c221obus));
wire [temp_w*7-1:0] c222ibus;
wire [data_w*7-1:0] c222obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU222 ( .en(en), .clk(clk), .rst(rst), .q(c222ibus), .r(c222obus));
wire [temp_w*7-1:0] c223ibus;
wire [data_w*7-1:0] c223obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU223 ( .en(en), .clk(clk), .rst(rst), .q(c223ibus), .r(c223obus));
wire [temp_w*7-1:0] c224ibus;
wire [data_w*7-1:0] c224obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU224 ( .en(en), .clk(clk), .rst(rst), .q(c224ibus), .r(c224obus));
wire [temp_w*7-1:0] c225ibus;
wire [data_w*7-1:0] c225obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU225 ( .en(en), .clk(clk), .rst(rst), .q(c225ibus), .r(c225obus));
wire [temp_w*7-1:0] c226ibus;
wire [data_w*7-1:0] c226obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU226 ( .en(en), .clk(clk), .rst(rst), .q(c226ibus), .r(c226obus));
wire [temp_w*7-1:0] c227ibus;
wire [data_w*7-1:0] c227obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU227 ( .en(en), .clk(clk), .rst(rst), .q(c227ibus), .r(c227obus));
wire [temp_w*7-1:0] c228ibus;
wire [data_w*7-1:0] c228obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU228 ( .en(en), .clk(clk), .rst(rst), .q(c228ibus), .r(c228obus));
wire [temp_w*7-1:0] c229ibus;
wire [data_w*7-1:0] c229obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU229 ( .en(en), .clk(clk), .rst(rst), .q(c229ibus), .r(c229obus));
wire [temp_w*7-1:0] c230ibus;
wire [data_w*7-1:0] c230obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU230 ( .en(en), .clk(clk), .rst(rst), .q(c230ibus), .r(c230obus));
wire [temp_w*7-1:0] c231ibus;
wire [data_w*7-1:0] c231obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU231 ( .en(en), .clk(clk), .rst(rst), .q(c231ibus), .r(c231obus));
wire [temp_w*7-1:0] c232ibus;
wire [data_w*7-1:0] c232obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU232 ( .en(en), .clk(clk), .rst(rst), .q(c232ibus), .r(c232obus));
wire [temp_w*7-1:0] c233ibus;
wire [data_w*7-1:0] c233obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU233 ( .en(en), .clk(clk), .rst(rst), .q(c233ibus), .r(c233obus));
wire [temp_w*7-1:0] c234ibus;
wire [data_w*7-1:0] c234obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU234 ( .en(en), .clk(clk), .rst(rst), .q(c234ibus), .r(c234obus));
wire [temp_w*7-1:0] c235ibus;
wire [data_w*7-1:0] c235obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU235 ( .en(en), .clk(clk), .rst(rst), .q(c235ibus), .r(c235obus));
wire [temp_w*7-1:0] c236ibus;
wire [data_w*7-1:0] c236obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU236 ( .en(en), .clk(clk), .rst(rst), .q(c236ibus), .r(c236obus));
wire [temp_w*7-1:0] c237ibus;
wire [data_w*7-1:0] c237obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU237 ( .en(en), .clk(clk), .rst(rst), .q(c237ibus), .r(c237obus));
wire [temp_w*7-1:0] c238ibus;
wire [data_w*7-1:0] c238obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU238 ( .en(en), .clk(clk), .rst(rst), .q(c238ibus), .r(c238obus));
wire [temp_w*7-1:0] c239ibus;
wire [data_w*7-1:0] c239obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU239 ( .en(en), .clk(clk), .rst(rst), .q(c239ibus), .r(c239obus));
wire [temp_w*7-1:0] c240ibus;
wire [data_w*7-1:0] c240obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU240 ( .en(en), .clk(clk), .rst(rst), .q(c240ibus), .r(c240obus));
wire [temp_w*7-1:0] c241ibus;
wire [data_w*7-1:0] c241obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU241 ( .en(en), .clk(clk), .rst(rst), .q(c241ibus), .r(c241obus));
wire [temp_w*7-1:0] c242ibus;
wire [data_w*7-1:0] c242obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU242 ( .en(en), .clk(clk), .rst(rst), .q(c242ibus), .r(c242obus));
wire [temp_w*7-1:0] c243ibus;
wire [data_w*7-1:0] c243obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU243 ( .en(en), .clk(clk), .rst(rst), .q(c243ibus), .r(c243obus));
wire [temp_w*7-1:0] c244ibus;
wire [data_w*7-1:0] c244obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU244 ( .en(en), .clk(clk), .rst(rst), .q(c244ibus), .r(c244obus));
wire [temp_w*7-1:0] c245ibus;
wire [data_w*7-1:0] c245obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU245 ( .en(en), .clk(clk), .rst(rst), .q(c245ibus), .r(c245obus));
wire [temp_w*7-1:0] c246ibus;
wire [data_w*7-1:0] c246obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU246 ( .en(en), .clk(clk), .rst(rst), .q(c246ibus), .r(c246obus));
wire [temp_w*7-1:0] c247ibus;
wire [data_w*7-1:0] c247obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU247 ( .en(en), .clk(clk), .rst(rst), .q(c247ibus), .r(c247obus));
wire [temp_w*7-1:0] c248ibus;
wire [data_w*7-1:0] c248obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU248 ( .en(en), .clk(clk), .rst(rst), .q(c248ibus), .r(c248obus));
wire [temp_w*7-1:0] c249ibus;
wire [data_w*7-1:0] c249obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU249 ( .en(en), .clk(clk), .rst(rst), .q(c249ibus), .r(c249obus));
wire [temp_w*7-1:0] c250ibus;
wire [data_w*7-1:0] c250obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU250 ( .en(en), .clk(clk), .rst(rst), .q(c250ibus), .r(c250obus));
wire [temp_w*7-1:0] c251ibus;
wire [data_w*7-1:0] c251obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU251 ( .en(en), .clk(clk), .rst(rst), .q(c251ibus), .r(c251obus));
wire [temp_w*7-1:0] c252ibus;
wire [data_w*7-1:0] c252obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU252 ( .en(en), .clk(clk), .rst(rst), .q(c252ibus), .r(c252obus));
wire [temp_w*7-1:0] c253ibus;
wire [data_w*7-1:0] c253obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU253 ( .en(en), .clk(clk), .rst(rst), .q(c253ibus), .r(c253obus));
wire [temp_w*7-1:0] c254ibus;
wire [data_w*7-1:0] c254obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU254 ( .en(en), .clk(clk), .rst(rst), .q(c254ibus), .r(c254obus));
wire [temp_w*7-1:0] c255ibus;
wire [data_w*7-1:0] c255obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU255 ( .en(en), .clk(clk), .rst(rst), .q(c255ibus), .r(c255obus));
wire [temp_w*7-1:0] c256ibus;
wire [data_w*7-1:0] c256obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU256 ( .en(en), .clk(clk), .rst(rst), .q(c256ibus), .r(c256obus));
wire [temp_w*7-1:0] c257ibus;
wire [data_w*7-1:0] c257obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU257 ( .en(en), .clk(clk), .rst(rst), .q(c257ibus), .r(c257obus));
wire [temp_w*7-1:0] c258ibus;
wire [data_w*7-1:0] c258obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU258 ( .en(en), .clk(clk), .rst(rst), .q(c258ibus), .r(c258obus));
wire [temp_w*7-1:0] c259ibus;
wire [data_w*7-1:0] c259obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU259 ( .en(en), .clk(clk), .rst(rst), .q(c259ibus), .r(c259obus));
wire [temp_w*7-1:0] c260ibus;
wire [data_w*7-1:0] c260obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU260 ( .en(en), .clk(clk), .rst(rst), .q(c260ibus), .r(c260obus));
wire [temp_w*7-1:0] c261ibus;
wire [data_w*7-1:0] c261obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU261 ( .en(en), .clk(clk), .rst(rst), .q(c261ibus), .r(c261obus));
wire [temp_w*7-1:0] c262ibus;
wire [data_w*7-1:0] c262obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU262 ( .en(en), .clk(clk), .rst(rst), .q(c262ibus), .r(c262obus));
wire [temp_w*7-1:0] c263ibus;
wire [data_w*7-1:0] c263obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU263 ( .en(en), .clk(clk), .rst(rst), .q(c263ibus), .r(c263obus));
wire [temp_w*7-1:0] c264ibus;
wire [data_w*7-1:0] c264obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU264 ( .en(en), .clk(clk), .rst(rst), .q(c264ibus), .r(c264obus));
wire [temp_w*7-1:0] c265ibus;
wire [data_w*7-1:0] c265obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU265 ( .en(en), .clk(clk), .rst(rst), .q(c265ibus), .r(c265obus));
wire [temp_w*7-1:0] c266ibus;
wire [data_w*7-1:0] c266obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU266 ( .en(en), .clk(clk), .rst(rst), .q(c266ibus), .r(c266obus));
wire [temp_w*7-1:0] c267ibus;
wire [data_w*7-1:0] c267obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU267 ( .en(en), .clk(clk), .rst(rst), .q(c267ibus), .r(c267obus));
wire [temp_w*7-1:0] c268ibus;
wire [data_w*7-1:0] c268obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU268 ( .en(en), .clk(clk), .rst(rst), .q(c268ibus), .r(c268obus));
wire [temp_w*7-1:0] c269ibus;
wire [data_w*7-1:0] c269obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU269 ( .en(en), .clk(clk), .rst(rst), .q(c269ibus), .r(c269obus));
wire [temp_w*7-1:0] c270ibus;
wire [data_w*7-1:0] c270obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU270 ( .en(en), .clk(clk), .rst(rst), .q(c270ibus), .r(c270obus));
wire [temp_w*7-1:0] c271ibus;
wire [data_w*7-1:0] c271obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU271 ( .en(en), .clk(clk), .rst(rst), .q(c271ibus), .r(c271obus));
wire [temp_w*7-1:0] c272ibus;
wire [data_w*7-1:0] c272obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU272 ( .en(en), .clk(clk), .rst(rst), .q(c272ibus), .r(c272obus));
wire [temp_w*7-1:0] c273ibus;
wire [data_w*7-1:0] c273obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU273 ( .en(en), .clk(clk), .rst(rst), .q(c273ibus), .r(c273obus));
wire [temp_w*7-1:0] c274ibus;
wire [data_w*7-1:0] c274obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU274 ( .en(en), .clk(clk), .rst(rst), .q(c274ibus), .r(c274obus));
wire [temp_w*7-1:0] c275ibus;
wire [data_w*7-1:0] c275obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU275 ( .en(en), .clk(clk), .rst(rst), .q(c275ibus), .r(c275obus));
wire [temp_w*7-1:0] c276ibus;
wire [data_w*7-1:0] c276obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU276 ( .en(en), .clk(clk), .rst(rst), .q(c276ibus), .r(c276obus));
wire [temp_w*7-1:0] c277ibus;
wire [data_w*7-1:0] c277obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU277 ( .en(en), .clk(clk), .rst(rst), .q(c277ibus), .r(c277obus));
wire [temp_w*7-1:0] c278ibus;
wire [data_w*7-1:0] c278obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU278 ( .en(en), .clk(clk), .rst(rst), .q(c278ibus), .r(c278obus));
wire [temp_w*7-1:0] c279ibus;
wire [data_w*7-1:0] c279obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU279 ( .en(en), .clk(clk), .rst(rst), .q(c279ibus), .r(c279obus));
wire [temp_w*7-1:0] c280ibus;
wire [data_w*7-1:0] c280obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU280 ( .en(en), .clk(clk), .rst(rst), .q(c280ibus), .r(c280obus));
wire [temp_w*7-1:0] c281ibus;
wire [data_w*7-1:0] c281obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU281 ( .en(en), .clk(clk), .rst(rst), .q(c281ibus), .r(c281obus));
wire [temp_w*7-1:0] c282ibus;
wire [data_w*7-1:0] c282obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU282 ( .en(en), .clk(clk), .rst(rst), .q(c282ibus), .r(c282obus));
wire [temp_w*7-1:0] c283ibus;
wire [data_w*7-1:0] c283obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU283 ( .en(en), .clk(clk), .rst(rst), .q(c283ibus), .r(c283obus));
wire [temp_w*7-1:0] c284ibus;
wire [data_w*7-1:0] c284obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU284 ( .en(en), .clk(clk), .rst(rst), .q(c284ibus), .r(c284obus));
wire [temp_w*7-1:0] c285ibus;
wire [data_w*7-1:0] c285obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU285 ( .en(en), .clk(clk), .rst(rst), .q(c285ibus), .r(c285obus));
wire [temp_w*7-1:0] c286ibus;
wire [data_w*7-1:0] c286obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU286 ( .en(en), .clk(clk), .rst(rst), .q(c286ibus), .r(c286obus));
wire [temp_w*7-1:0] c287ibus;
wire [data_w*7-1:0] c287obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU287 ( .en(en), .clk(clk), .rst(rst), .q(c287ibus), .r(c287obus));
wire [temp_w*6-1:0] c288ibus;
wire [data_w*6-1:0] c288obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU288 ( .en(en), .clk(clk), .rst(rst), .q(c288ibus), .r(c288obus));
wire [temp_w*6-1:0] c289ibus;
wire [data_w*6-1:0] c289obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU289 ( .en(en), .clk(clk), .rst(rst), .q(c289ibus), .r(c289obus));
wire [temp_w*6-1:0] c290ibus;
wire [data_w*6-1:0] c290obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU290 ( .en(en), .clk(clk), .rst(rst), .q(c290ibus), .r(c290obus));
wire [temp_w*6-1:0] c291ibus;
wire [data_w*6-1:0] c291obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU291 ( .en(en), .clk(clk), .rst(rst), .q(c291ibus), .r(c291obus));
wire [temp_w*6-1:0] c292ibus;
wire [data_w*6-1:0] c292obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU292 ( .en(en), .clk(clk), .rst(rst), .q(c292ibus), .r(c292obus));
wire [temp_w*6-1:0] c293ibus;
wire [data_w*6-1:0] c293obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU293 ( .en(en), .clk(clk), .rst(rst), .q(c293ibus), .r(c293obus));
wire [temp_w*6-1:0] c294ibus;
wire [data_w*6-1:0] c294obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU294 ( .en(en), .clk(clk), .rst(rst), .q(c294ibus), .r(c294obus));
wire [temp_w*6-1:0] c295ibus;
wire [data_w*6-1:0] c295obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU295 ( .en(en), .clk(clk), .rst(rst), .q(c295ibus), .r(c295obus));
wire [temp_w*6-1:0] c296ibus;
wire [data_w*6-1:0] c296obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU296 ( .en(en), .clk(clk), .rst(rst), .q(c296ibus), .r(c296obus));
wire [temp_w*6-1:0] c297ibus;
wire [data_w*6-1:0] c297obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU297 ( .en(en), .clk(clk), .rst(rst), .q(c297ibus), .r(c297obus));
wire [temp_w*6-1:0] c298ibus;
wire [data_w*6-1:0] c298obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU298 ( .en(en), .clk(clk), .rst(rst), .q(c298ibus), .r(c298obus));
wire [temp_w*6-1:0] c299ibus;
wire [data_w*6-1:0] c299obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU299 ( .en(en), .clk(clk), .rst(rst), .q(c299ibus), .r(c299obus));
wire [temp_w*6-1:0] c300ibus;
wire [data_w*6-1:0] c300obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU300 ( .en(en), .clk(clk), .rst(rst), .q(c300ibus), .r(c300obus));
wire [temp_w*6-1:0] c301ibus;
wire [data_w*6-1:0] c301obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU301 ( .en(en), .clk(clk), .rst(rst), .q(c301ibus), .r(c301obus));
wire [temp_w*6-1:0] c302ibus;
wire [data_w*6-1:0] c302obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU302 ( .en(en), .clk(clk), .rst(rst), .q(c302ibus), .r(c302obus));
wire [temp_w*6-1:0] c303ibus;
wire [data_w*6-1:0] c303obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU303 ( .en(en), .clk(clk), .rst(rst), .q(c303ibus), .r(c303obus));
wire [temp_w*6-1:0] c304ibus;
wire [data_w*6-1:0] c304obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU304 ( .en(en), .clk(clk), .rst(rst), .q(c304ibus), .r(c304obus));
wire [temp_w*6-1:0] c305ibus;
wire [data_w*6-1:0] c305obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU305 ( .en(en), .clk(clk), .rst(rst), .q(c305ibus), .r(c305obus));
wire [temp_w*6-1:0] c306ibus;
wire [data_w*6-1:0] c306obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU306 ( .en(en), .clk(clk), .rst(rst), .q(c306ibus), .r(c306obus));
wire [temp_w*6-1:0] c307ibus;
wire [data_w*6-1:0] c307obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU307 ( .en(en), .clk(clk), .rst(rst), .q(c307ibus), .r(c307obus));
wire [temp_w*6-1:0] c308ibus;
wire [data_w*6-1:0] c308obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU308 ( .en(en), .clk(clk), .rst(rst), .q(c308ibus), .r(c308obus));
wire [temp_w*6-1:0] c309ibus;
wire [data_w*6-1:0] c309obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU309 ( .en(en), .clk(clk), .rst(rst), .q(c309ibus), .r(c309obus));
wire [temp_w*6-1:0] c310ibus;
wire [data_w*6-1:0] c310obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU310 ( .en(en), .clk(clk), .rst(rst), .q(c310ibus), .r(c310obus));
wire [temp_w*6-1:0] c311ibus;
wire [data_w*6-1:0] c311obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU311 ( .en(en), .clk(clk), .rst(rst), .q(c311ibus), .r(c311obus));
wire [temp_w*6-1:0] c312ibus;
wire [data_w*6-1:0] c312obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU312 ( .en(en), .clk(clk), .rst(rst), .q(c312ibus), .r(c312obus));
wire [temp_w*6-1:0] c313ibus;
wire [data_w*6-1:0] c313obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU313 ( .en(en), .clk(clk), .rst(rst), .q(c313ibus), .r(c313obus));
wire [temp_w*6-1:0] c314ibus;
wire [data_w*6-1:0] c314obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU314 ( .en(en), .clk(clk), .rst(rst), .q(c314ibus), .r(c314obus));
wire [temp_w*6-1:0] c315ibus;
wire [data_w*6-1:0] c315obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU315 ( .en(en), .clk(clk), .rst(rst), .q(c315ibus), .r(c315obus));
wire [temp_w*6-1:0] c316ibus;
wire [data_w*6-1:0] c316obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU316 ( .en(en), .clk(clk), .rst(rst), .q(c316ibus), .r(c316obus));
wire [temp_w*6-1:0] c317ibus;
wire [data_w*6-1:0] c317obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU317 ( .en(en), .clk(clk), .rst(rst), .q(c317ibus), .r(c317obus));
wire [temp_w*6-1:0] c318ibus;
wire [data_w*6-1:0] c318obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU318 ( .en(en), .clk(clk), .rst(rst), .q(c318ibus), .r(c318obus));
wire [temp_w*6-1:0] c319ibus;
wire [data_w*6-1:0] c319obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU319 ( .en(en), .clk(clk), .rst(rst), .q(c319ibus), .r(c319obus));
wire [temp_w*6-1:0] c320ibus;
wire [data_w*6-1:0] c320obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU320 ( .en(en), .clk(clk), .rst(rst), .q(c320ibus), .r(c320obus));
wire [temp_w*6-1:0] c321ibus;
wire [data_w*6-1:0] c321obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU321 ( .en(en), .clk(clk), .rst(rst), .q(c321ibus), .r(c321obus));
wire [temp_w*6-1:0] c322ibus;
wire [data_w*6-1:0] c322obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU322 ( .en(en), .clk(clk), .rst(rst), .q(c322ibus), .r(c322obus));
wire [temp_w*6-1:0] c323ibus;
wire [data_w*6-1:0] c323obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU323 ( .en(en), .clk(clk), .rst(rst), .q(c323ibus), .r(c323obus));
wire [temp_w*6-1:0] c324ibus;
wire [data_w*6-1:0] c324obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU324 ( .en(en), .clk(clk), .rst(rst), .q(c324ibus), .r(c324obus));
wire [temp_w*6-1:0] c325ibus;
wire [data_w*6-1:0] c325obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU325 ( .en(en), .clk(clk), .rst(rst), .q(c325ibus), .r(c325obus));
wire [temp_w*6-1:0] c326ibus;
wire [data_w*6-1:0] c326obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU326 ( .en(en), .clk(clk), .rst(rst), .q(c326ibus), .r(c326obus));
wire [temp_w*6-1:0] c327ibus;
wire [data_w*6-1:0] c327obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU327 ( .en(en), .clk(clk), .rst(rst), .q(c327ibus), .r(c327obus));
wire [temp_w*6-1:0] c328ibus;
wire [data_w*6-1:0] c328obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU328 ( .en(en), .clk(clk), .rst(rst), .q(c328ibus), .r(c328obus));
wire [temp_w*6-1:0] c329ibus;
wire [data_w*6-1:0] c329obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU329 ( .en(en), .clk(clk), .rst(rst), .q(c329ibus), .r(c329obus));
wire [temp_w*6-1:0] c330ibus;
wire [data_w*6-1:0] c330obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU330 ( .en(en), .clk(clk), .rst(rst), .q(c330ibus), .r(c330obus));
wire [temp_w*6-1:0] c331ibus;
wire [data_w*6-1:0] c331obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU331 ( .en(en), .clk(clk), .rst(rst), .q(c331ibus), .r(c331obus));
wire [temp_w*6-1:0] c332ibus;
wire [data_w*6-1:0] c332obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU332 ( .en(en), .clk(clk), .rst(rst), .q(c332ibus), .r(c332obus));
wire [temp_w*6-1:0] c333ibus;
wire [data_w*6-1:0] c333obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU333 ( .en(en), .clk(clk), .rst(rst), .q(c333ibus), .r(c333obus));
wire [temp_w*6-1:0] c334ibus;
wire [data_w*6-1:0] c334obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU334 ( .en(en), .clk(clk), .rst(rst), .q(c334ibus), .r(c334obus));
wire [temp_w*6-1:0] c335ibus;
wire [data_w*6-1:0] c335obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU335 ( .en(en), .clk(clk), .rst(rst), .q(c335ibus), .r(c335obus));
wire [temp_w*6-1:0] c336ibus;
wire [data_w*6-1:0] c336obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU336 ( .en(en), .clk(clk), .rst(rst), .q(c336ibus), .r(c336obus));
wire [temp_w*6-1:0] c337ibus;
wire [data_w*6-1:0] c337obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU337 ( .en(en), .clk(clk), .rst(rst), .q(c337ibus), .r(c337obus));
wire [temp_w*6-1:0] c338ibus;
wire [data_w*6-1:0] c338obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU338 ( .en(en), .clk(clk), .rst(rst), .q(c338ibus), .r(c338obus));
wire [temp_w*6-1:0] c339ibus;
wire [data_w*6-1:0] c339obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU339 ( .en(en), .clk(clk), .rst(rst), .q(c339ibus), .r(c339obus));
wire [temp_w*6-1:0] c340ibus;
wire [data_w*6-1:0] c340obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU340 ( .en(en), .clk(clk), .rst(rst), .q(c340ibus), .r(c340obus));
wire [temp_w*6-1:0] c341ibus;
wire [data_w*6-1:0] c341obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU341 ( .en(en), .clk(clk), .rst(rst), .q(c341ibus), .r(c341obus));
wire [temp_w*6-1:0] c342ibus;
wire [data_w*6-1:0] c342obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU342 ( .en(en), .clk(clk), .rst(rst), .q(c342ibus), .r(c342obus));
wire [temp_w*6-1:0] c343ibus;
wire [data_w*6-1:0] c343obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU343 ( .en(en), .clk(clk), .rst(rst), .q(c343ibus), .r(c343obus));
wire [temp_w*6-1:0] c344ibus;
wire [data_w*6-1:0] c344obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU344 ( .en(en), .clk(clk), .rst(rst), .q(c344ibus), .r(c344obus));
wire [temp_w*6-1:0] c345ibus;
wire [data_w*6-1:0] c345obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU345 ( .en(en), .clk(clk), .rst(rst), .q(c345ibus), .r(c345obus));
wire [temp_w*6-1:0] c346ibus;
wire [data_w*6-1:0] c346obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU346 ( .en(en), .clk(clk), .rst(rst), .q(c346ibus), .r(c346obus));
wire [temp_w*6-1:0] c347ibus;
wire [data_w*6-1:0] c347obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU347 ( .en(en), .clk(clk), .rst(rst), .q(c347ibus), .r(c347obus));
wire [temp_w*6-1:0] c348ibus;
wire [data_w*6-1:0] c348obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU348 ( .en(en), .clk(clk), .rst(rst), .q(c348ibus), .r(c348obus));
wire [temp_w*6-1:0] c349ibus;
wire [data_w*6-1:0] c349obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU349 ( .en(en), .clk(clk), .rst(rst), .q(c349ibus), .r(c349obus));
wire [temp_w*6-1:0] c350ibus;
wire [data_w*6-1:0] c350obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU350 ( .en(en), .clk(clk), .rst(rst), .q(c350ibus), .r(c350obus));
wire [temp_w*6-1:0] c351ibus;
wire [data_w*6-1:0] c351obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU351 ( .en(en), .clk(clk), .rst(rst), .q(c351ibus), .r(c351obus));
wire [temp_w*6-1:0] c352ibus;
wire [data_w*6-1:0] c352obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU352 ( .en(en), .clk(clk), .rst(rst), .q(c352ibus), .r(c352obus));
wire [temp_w*6-1:0] c353ibus;
wire [data_w*6-1:0] c353obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU353 ( .en(en), .clk(clk), .rst(rst), .q(c353ibus), .r(c353obus));
wire [temp_w*6-1:0] c354ibus;
wire [data_w*6-1:0] c354obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU354 ( .en(en), .clk(clk), .rst(rst), .q(c354ibus), .r(c354obus));
wire [temp_w*6-1:0] c355ibus;
wire [data_w*6-1:0] c355obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU355 ( .en(en), .clk(clk), .rst(rst), .q(c355ibus), .r(c355obus));
wire [temp_w*6-1:0] c356ibus;
wire [data_w*6-1:0] c356obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU356 ( .en(en), .clk(clk), .rst(rst), .q(c356ibus), .r(c356obus));
wire [temp_w*6-1:0] c357ibus;
wire [data_w*6-1:0] c357obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU357 ( .en(en), .clk(clk), .rst(rst), .q(c357ibus), .r(c357obus));
wire [temp_w*6-1:0] c358ibus;
wire [data_w*6-1:0] c358obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU358 ( .en(en), .clk(clk), .rst(rst), .q(c358ibus), .r(c358obus));
wire [temp_w*6-1:0] c359ibus;
wire [data_w*6-1:0] c359obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU359 ( .en(en), .clk(clk), .rst(rst), .q(c359ibus), .r(c359obus));
wire [temp_w*6-1:0] c360ibus;
wire [data_w*6-1:0] c360obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU360 ( .en(en), .clk(clk), .rst(rst), .q(c360ibus), .r(c360obus));
wire [temp_w*6-1:0] c361ibus;
wire [data_w*6-1:0] c361obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU361 ( .en(en), .clk(clk), .rst(rst), .q(c361ibus), .r(c361obus));
wire [temp_w*6-1:0] c362ibus;
wire [data_w*6-1:0] c362obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU362 ( .en(en), .clk(clk), .rst(rst), .q(c362ibus), .r(c362obus));
wire [temp_w*6-1:0] c363ibus;
wire [data_w*6-1:0] c363obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU363 ( .en(en), .clk(clk), .rst(rst), .q(c363ibus), .r(c363obus));
wire [temp_w*6-1:0] c364ibus;
wire [data_w*6-1:0] c364obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU364 ( .en(en), .clk(clk), .rst(rst), .q(c364ibus), .r(c364obus));
wire [temp_w*6-1:0] c365ibus;
wire [data_w*6-1:0] c365obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU365 ( .en(en), .clk(clk), .rst(rst), .q(c365ibus), .r(c365obus));
wire [temp_w*6-1:0] c366ibus;
wire [data_w*6-1:0] c366obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU366 ( .en(en), .clk(clk), .rst(rst), .q(c366ibus), .r(c366obus));
wire [temp_w*6-1:0] c367ibus;
wire [data_w*6-1:0] c367obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU367 ( .en(en), .clk(clk), .rst(rst), .q(c367ibus), .r(c367obus));
wire [temp_w*6-1:0] c368ibus;
wire [data_w*6-1:0] c368obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU368 ( .en(en), .clk(clk), .rst(rst), .q(c368ibus), .r(c368obus));
wire [temp_w*6-1:0] c369ibus;
wire [data_w*6-1:0] c369obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU369 ( .en(en), .clk(clk), .rst(rst), .q(c369ibus), .r(c369obus));
wire [temp_w*6-1:0] c370ibus;
wire [data_w*6-1:0] c370obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU370 ( .en(en), .clk(clk), .rst(rst), .q(c370ibus), .r(c370obus));
wire [temp_w*6-1:0] c371ibus;
wire [data_w*6-1:0] c371obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU371 ( .en(en), .clk(clk), .rst(rst), .q(c371ibus), .r(c371obus));
wire [temp_w*6-1:0] c372ibus;
wire [data_w*6-1:0] c372obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU372 ( .en(en), .clk(clk), .rst(rst), .q(c372ibus), .r(c372obus));
wire [temp_w*6-1:0] c373ibus;
wire [data_w*6-1:0] c373obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU373 ( .en(en), .clk(clk), .rst(rst), .q(c373ibus), .r(c373obus));
wire [temp_w*6-1:0] c374ibus;
wire [data_w*6-1:0] c374obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU374 ( .en(en), .clk(clk), .rst(rst), .q(c374ibus), .r(c374obus));
wire [temp_w*6-1:0] c375ibus;
wire [data_w*6-1:0] c375obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU375 ( .en(en), .clk(clk), .rst(rst), .q(c375ibus), .r(c375obus));
wire [temp_w*6-1:0] c376ibus;
wire [data_w*6-1:0] c376obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU376 ( .en(en), .clk(clk), .rst(rst), .q(c376ibus), .r(c376obus));
wire [temp_w*6-1:0] c377ibus;
wire [data_w*6-1:0] c377obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU377 ( .en(en), .clk(clk), .rst(rst), .q(c377ibus), .r(c377obus));
wire [temp_w*6-1:0] c378ibus;
wire [data_w*6-1:0] c378obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU378 ( .en(en), .clk(clk), .rst(rst), .q(c378ibus), .r(c378obus));
wire [temp_w*6-1:0] c379ibus;
wire [data_w*6-1:0] c379obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU379 ( .en(en), .clk(clk), .rst(rst), .q(c379ibus), .r(c379obus));
wire [temp_w*6-1:0] c380ibus;
wire [data_w*6-1:0] c380obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU380 ( .en(en), .clk(clk), .rst(rst), .q(c380ibus), .r(c380obus));
wire [temp_w*6-1:0] c381ibus;
wire [data_w*6-1:0] c381obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU381 ( .en(en), .clk(clk), .rst(rst), .q(c381ibus), .r(c381obus));
wire [temp_w*6-1:0] c382ibus;
wire [data_w*6-1:0] c382obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU382 ( .en(en), .clk(clk), .rst(rst), .q(c382ibus), .r(c382obus));
wire [temp_w*6-1:0] c383ibus;
wire [data_w*6-1:0] c383obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU383 ( .en(en), .clk(clk), .rst(rst), .q(c383ibus), .r(c383obus));
wire [temp_w*6-1:0] c384ibus;
wire [data_w*6-1:0] c384obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU384 ( .en(en), .clk(clk), .rst(rst), .q(c384ibus), .r(c384obus));
wire [temp_w*6-1:0] c385ibus;
wire [data_w*6-1:0] c385obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU385 ( .en(en), .clk(clk), .rst(rst), .q(c385ibus), .r(c385obus));
wire [temp_w*6-1:0] c386ibus;
wire [data_w*6-1:0] c386obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU386 ( .en(en), .clk(clk), .rst(rst), .q(c386ibus), .r(c386obus));
wire [temp_w*6-1:0] c387ibus;
wire [data_w*6-1:0] c387obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU387 ( .en(en), .clk(clk), .rst(rst), .q(c387ibus), .r(c387obus));
wire [temp_w*6-1:0] c388ibus;
wire [data_w*6-1:0] c388obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU388 ( .en(en), .clk(clk), .rst(rst), .q(c388ibus), .r(c388obus));
wire [temp_w*6-1:0] c389ibus;
wire [data_w*6-1:0] c389obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU389 ( .en(en), .clk(clk), .rst(rst), .q(c389ibus), .r(c389obus));
wire [temp_w*6-1:0] c390ibus;
wire [data_w*6-1:0] c390obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU390 ( .en(en), .clk(clk), .rst(rst), .q(c390ibus), .r(c390obus));
wire [temp_w*6-1:0] c391ibus;
wire [data_w*6-1:0] c391obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU391 ( .en(en), .clk(clk), .rst(rst), .q(c391ibus), .r(c391obus));
wire [temp_w*6-1:0] c392ibus;
wire [data_w*6-1:0] c392obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU392 ( .en(en), .clk(clk), .rst(rst), .q(c392ibus), .r(c392obus));
wire [temp_w*6-1:0] c393ibus;
wire [data_w*6-1:0] c393obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU393 ( .en(en), .clk(clk), .rst(rst), .q(c393ibus), .r(c393obus));
wire [temp_w*6-1:0] c394ibus;
wire [data_w*6-1:0] c394obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU394 ( .en(en), .clk(clk), .rst(rst), .q(c394ibus), .r(c394obus));
wire [temp_w*6-1:0] c395ibus;
wire [data_w*6-1:0] c395obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU395 ( .en(en), .clk(clk), .rst(rst), .q(c395ibus), .r(c395obus));
wire [temp_w*6-1:0] c396ibus;
wire [data_w*6-1:0] c396obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU396 ( .en(en), .clk(clk), .rst(rst), .q(c396ibus), .r(c396obus));
wire [temp_w*6-1:0] c397ibus;
wire [data_w*6-1:0] c397obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU397 ( .en(en), .clk(clk), .rst(rst), .q(c397ibus), .r(c397obus));
wire [temp_w*6-1:0] c398ibus;
wire [data_w*6-1:0] c398obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU398 ( .en(en), .clk(clk), .rst(rst), .q(c398ibus), .r(c398obus));
wire [temp_w*6-1:0] c399ibus;
wire [data_w*6-1:0] c399obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU399 ( .en(en), .clk(clk), .rst(rst), .q(c399ibus), .r(c399obus));
wire [temp_w*6-1:0] c400ibus;
wire [data_w*6-1:0] c400obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU400 ( .en(en), .clk(clk), .rst(rst), .q(c400ibus), .r(c400obus));
wire [temp_w*6-1:0] c401ibus;
wire [data_w*6-1:0] c401obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU401 ( .en(en), .clk(clk), .rst(rst), .q(c401ibus), .r(c401obus));
wire [temp_w*6-1:0] c402ibus;
wire [data_w*6-1:0] c402obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU402 ( .en(en), .clk(clk), .rst(rst), .q(c402ibus), .r(c402obus));
wire [temp_w*6-1:0] c403ibus;
wire [data_w*6-1:0] c403obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU403 ( .en(en), .clk(clk), .rst(rst), .q(c403ibus), .r(c403obus));
wire [temp_w*6-1:0] c404ibus;
wire [data_w*6-1:0] c404obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU404 ( .en(en), .clk(clk), .rst(rst), .q(c404ibus), .r(c404obus));
wire [temp_w*6-1:0] c405ibus;
wire [data_w*6-1:0] c405obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU405 ( .en(en), .clk(clk), .rst(rst), .q(c405ibus), .r(c405obus));
wire [temp_w*6-1:0] c406ibus;
wire [data_w*6-1:0] c406obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU406 ( .en(en), .clk(clk), .rst(rst), .q(c406ibus), .r(c406obus));
wire [temp_w*6-1:0] c407ibus;
wire [data_w*6-1:0] c407obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU407 ( .en(en), .clk(clk), .rst(rst), .q(c407ibus), .r(c407obus));
wire [temp_w*6-1:0] c408ibus;
wire [data_w*6-1:0] c408obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU408 ( .en(en), .clk(clk), .rst(rst), .q(c408ibus), .r(c408obus));
wire [temp_w*6-1:0] c409ibus;
wire [data_w*6-1:0] c409obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU409 ( .en(en), .clk(clk), .rst(rst), .q(c409ibus), .r(c409obus));
wire [temp_w*6-1:0] c410ibus;
wire [data_w*6-1:0] c410obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU410 ( .en(en), .clk(clk), .rst(rst), .q(c410ibus), .r(c410obus));
wire [temp_w*6-1:0] c411ibus;
wire [data_w*6-1:0] c411obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU411 ( .en(en), .clk(clk), .rst(rst), .q(c411ibus), .r(c411obus));
wire [temp_w*6-1:0] c412ibus;
wire [data_w*6-1:0] c412obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU412 ( .en(en), .clk(clk), .rst(rst), .q(c412ibus), .r(c412obus));
wire [temp_w*6-1:0] c413ibus;
wire [data_w*6-1:0] c413obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU413 ( .en(en), .clk(clk), .rst(rst), .q(c413ibus), .r(c413obus));
wire [temp_w*6-1:0] c414ibus;
wire [data_w*6-1:0] c414obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU414 ( .en(en), .clk(clk), .rst(rst), .q(c414ibus), .r(c414obus));
wire [temp_w*6-1:0] c415ibus;
wire [data_w*6-1:0] c415obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU415 ( .en(en), .clk(clk), .rst(rst), .q(c415ibus), .r(c415obus));
wire [temp_w*6-1:0] c416ibus;
wire [data_w*6-1:0] c416obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU416 ( .en(en), .clk(clk), .rst(rst), .q(c416ibus), .r(c416obus));
wire [temp_w*6-1:0] c417ibus;
wire [data_w*6-1:0] c417obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU417 ( .en(en), .clk(clk), .rst(rst), .q(c417ibus), .r(c417obus));
wire [temp_w*6-1:0] c418ibus;
wire [data_w*6-1:0] c418obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU418 ( .en(en), .clk(clk), .rst(rst), .q(c418ibus), .r(c418obus));
wire [temp_w*6-1:0] c419ibus;
wire [data_w*6-1:0] c419obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU419 ( .en(en), .clk(clk), .rst(rst), .q(c419ibus), .r(c419obus));
wire [temp_w*6-1:0] c420ibus;
wire [data_w*6-1:0] c420obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU420 ( .en(en), .clk(clk), .rst(rst), .q(c420ibus), .r(c420obus));
wire [temp_w*6-1:0] c421ibus;
wire [data_w*6-1:0] c421obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU421 ( .en(en), .clk(clk), .rst(rst), .q(c421ibus), .r(c421obus));
wire [temp_w*6-1:0] c422ibus;
wire [data_w*6-1:0] c422obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU422 ( .en(en), .clk(clk), .rst(rst), .q(c422ibus), .r(c422obus));
wire [temp_w*6-1:0] c423ibus;
wire [data_w*6-1:0] c423obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU423 ( .en(en), .clk(clk), .rst(rst), .q(c423ibus), .r(c423obus));
wire [temp_w*6-1:0] c424ibus;
wire [data_w*6-1:0] c424obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU424 ( .en(en), .clk(clk), .rst(rst), .q(c424ibus), .r(c424obus));
wire [temp_w*6-1:0] c425ibus;
wire [data_w*6-1:0] c425obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU425 ( .en(en), .clk(clk), .rst(rst), .q(c425ibus), .r(c425obus));
wire [temp_w*6-1:0] c426ibus;
wire [data_w*6-1:0] c426obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU426 ( .en(en), .clk(clk), .rst(rst), .q(c426ibus), .r(c426obus));
wire [temp_w*6-1:0] c427ibus;
wire [data_w*6-1:0] c427obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU427 ( .en(en), .clk(clk), .rst(rst), .q(c427ibus), .r(c427obus));
wire [temp_w*6-1:0] c428ibus;
wire [data_w*6-1:0] c428obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU428 ( .en(en), .clk(clk), .rst(rst), .q(c428ibus), .r(c428obus));
wire [temp_w*6-1:0] c429ibus;
wire [data_w*6-1:0] c429obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU429 ( .en(en), .clk(clk), .rst(rst), .q(c429ibus), .r(c429obus));
wire [temp_w*6-1:0] c430ibus;
wire [data_w*6-1:0] c430obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU430 ( .en(en), .clk(clk), .rst(rst), .q(c430ibus), .r(c430obus));
wire [temp_w*6-1:0] c431ibus;
wire [data_w*6-1:0] c431obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU431 ( .en(en), .clk(clk), .rst(rst), .q(c431ibus), .r(c431obus));
wire [temp_w*6-1:0] c432ibus;
wire [data_w*6-1:0] c432obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU432 ( .en(en), .clk(clk), .rst(rst), .q(c432ibus), .r(c432obus));
wire [temp_w*6-1:0] c433ibus;
wire [data_w*6-1:0] c433obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU433 ( .en(en), .clk(clk), .rst(rst), .q(c433ibus), .r(c433obus));
wire [temp_w*6-1:0] c434ibus;
wire [data_w*6-1:0] c434obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU434 ( .en(en), .clk(clk), .rst(rst), .q(c434ibus), .r(c434obus));
wire [temp_w*6-1:0] c435ibus;
wire [data_w*6-1:0] c435obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU435 ( .en(en), .clk(clk), .rst(rst), .q(c435ibus), .r(c435obus));
wire [temp_w*6-1:0] c436ibus;
wire [data_w*6-1:0] c436obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU436 ( .en(en), .clk(clk), .rst(rst), .q(c436ibus), .r(c436obus));
wire [temp_w*6-1:0] c437ibus;
wire [data_w*6-1:0] c437obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU437 ( .en(en), .clk(clk), .rst(rst), .q(c437ibus), .r(c437obus));
wire [temp_w*6-1:0] c438ibus;
wire [data_w*6-1:0] c438obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU438 ( .en(en), .clk(clk), .rst(rst), .q(c438ibus), .r(c438obus));
wire [temp_w*6-1:0] c439ibus;
wire [data_w*6-1:0] c439obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU439 ( .en(en), .clk(clk), .rst(rst), .q(c439ibus), .r(c439obus));
wire [temp_w*6-1:0] c440ibus;
wire [data_w*6-1:0] c440obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU440 ( .en(en), .clk(clk), .rst(rst), .q(c440ibus), .r(c440obus));
wire [temp_w*6-1:0] c441ibus;
wire [data_w*6-1:0] c441obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU441 ( .en(en), .clk(clk), .rst(rst), .q(c441ibus), .r(c441obus));
wire [temp_w*6-1:0] c442ibus;
wire [data_w*6-1:0] c442obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU442 ( .en(en), .clk(clk), .rst(rst), .q(c442ibus), .r(c442obus));
wire [temp_w*6-1:0] c443ibus;
wire [data_w*6-1:0] c443obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU443 ( .en(en), .clk(clk), .rst(rst), .q(c443ibus), .r(c443obus));
wire [temp_w*6-1:0] c444ibus;
wire [data_w*6-1:0] c444obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU444 ( .en(en), .clk(clk), .rst(rst), .q(c444ibus), .r(c444obus));
wire [temp_w*6-1:0] c445ibus;
wire [data_w*6-1:0] c445obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU445 ( .en(en), .clk(clk), .rst(rst), .q(c445ibus), .r(c445obus));
wire [temp_w*6-1:0] c446ibus;
wire [data_w*6-1:0] c446obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU446 ( .en(en), .clk(clk), .rst(rst), .q(c446ibus), .r(c446obus));
wire [temp_w*6-1:0] c447ibus;
wire [data_w*6-1:0] c447obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU447 ( .en(en), .clk(clk), .rst(rst), .q(c447ibus), .r(c447obus));
wire [temp_w*6-1:0] c448ibus;
wire [data_w*6-1:0] c448obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU448 ( .en(en), .clk(clk), .rst(rst), .q(c448ibus), .r(c448obus));
wire [temp_w*6-1:0] c449ibus;
wire [data_w*6-1:0] c449obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU449 ( .en(en), .clk(clk), .rst(rst), .q(c449ibus), .r(c449obus));
wire [temp_w*6-1:0] c450ibus;
wire [data_w*6-1:0] c450obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU450 ( .en(en), .clk(clk), .rst(rst), .q(c450ibus), .r(c450obus));
wire [temp_w*6-1:0] c451ibus;
wire [data_w*6-1:0] c451obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU451 ( .en(en), .clk(clk), .rst(rst), .q(c451ibus), .r(c451obus));
wire [temp_w*6-1:0] c452ibus;
wire [data_w*6-1:0] c452obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU452 ( .en(en), .clk(clk), .rst(rst), .q(c452ibus), .r(c452obus));
wire [temp_w*6-1:0] c453ibus;
wire [data_w*6-1:0] c453obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU453 ( .en(en), .clk(clk), .rst(rst), .q(c453ibus), .r(c453obus));
wire [temp_w*6-1:0] c454ibus;
wire [data_w*6-1:0] c454obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU454 ( .en(en), .clk(clk), .rst(rst), .q(c454ibus), .r(c454obus));
wire [temp_w*6-1:0] c455ibus;
wire [data_w*6-1:0] c455obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU455 ( .en(en), .clk(clk), .rst(rst), .q(c455ibus), .r(c455obus));
wire [temp_w*6-1:0] c456ibus;
wire [data_w*6-1:0] c456obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU456 ( .en(en), .clk(clk), .rst(rst), .q(c456ibus), .r(c456obus));
wire [temp_w*6-1:0] c457ibus;
wire [data_w*6-1:0] c457obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU457 ( .en(en), .clk(clk), .rst(rst), .q(c457ibus), .r(c457obus));
wire [temp_w*6-1:0] c458ibus;
wire [data_w*6-1:0] c458obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU458 ( .en(en), .clk(clk), .rst(rst), .q(c458ibus), .r(c458obus));
wire [temp_w*6-1:0] c459ibus;
wire [data_w*6-1:0] c459obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU459 ( .en(en), .clk(clk), .rst(rst), .q(c459ibus), .r(c459obus));
wire [temp_w*6-1:0] c460ibus;
wire [data_w*6-1:0] c460obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU460 ( .en(en), .clk(clk), .rst(rst), .q(c460ibus), .r(c460obus));
wire [temp_w*6-1:0] c461ibus;
wire [data_w*6-1:0] c461obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU461 ( .en(en), .clk(clk), .rst(rst), .q(c461ibus), .r(c461obus));
wire [temp_w*6-1:0] c462ibus;
wire [data_w*6-1:0] c462obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU462 ( .en(en), .clk(clk), .rst(rst), .q(c462ibus), .r(c462obus));
wire [temp_w*6-1:0] c463ibus;
wire [data_w*6-1:0] c463obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU463 ( .en(en), .clk(clk), .rst(rst), .q(c463ibus), .r(c463obus));
wire [temp_w*6-1:0] c464ibus;
wire [data_w*6-1:0] c464obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU464 ( .en(en), .clk(clk), .rst(rst), .q(c464ibus), .r(c464obus));
wire [temp_w*6-1:0] c465ibus;
wire [data_w*6-1:0] c465obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU465 ( .en(en), .clk(clk), .rst(rst), .q(c465ibus), .r(c465obus));
wire [temp_w*6-1:0] c466ibus;
wire [data_w*6-1:0] c466obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU466 ( .en(en), .clk(clk), .rst(rst), .q(c466ibus), .r(c466obus));
wire [temp_w*6-1:0] c467ibus;
wire [data_w*6-1:0] c467obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU467 ( .en(en), .clk(clk), .rst(rst), .q(c467ibus), .r(c467obus));
wire [temp_w*6-1:0] c468ibus;
wire [data_w*6-1:0] c468obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU468 ( .en(en), .clk(clk), .rst(rst), .q(c468ibus), .r(c468obus));
wire [temp_w*6-1:0] c469ibus;
wire [data_w*6-1:0] c469obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU469 ( .en(en), .clk(clk), .rst(rst), .q(c469ibus), .r(c469obus));
wire [temp_w*6-1:0] c470ibus;
wire [data_w*6-1:0] c470obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU470 ( .en(en), .clk(clk), .rst(rst), .q(c470ibus), .r(c470obus));
wire [temp_w*6-1:0] c471ibus;
wire [data_w*6-1:0] c471obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU471 ( .en(en), .clk(clk), .rst(rst), .q(c471ibus), .r(c471obus));
wire [temp_w*6-1:0] c472ibus;
wire [data_w*6-1:0] c472obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU472 ( .en(en), .clk(clk), .rst(rst), .q(c472ibus), .r(c472obus));
wire [temp_w*6-1:0] c473ibus;
wire [data_w*6-1:0] c473obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU473 ( .en(en), .clk(clk), .rst(rst), .q(c473ibus), .r(c473obus));
wire [temp_w*6-1:0] c474ibus;
wire [data_w*6-1:0] c474obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU474 ( .en(en), .clk(clk), .rst(rst), .q(c474ibus), .r(c474obus));
wire [temp_w*6-1:0] c475ibus;
wire [data_w*6-1:0] c475obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU475 ( .en(en), .clk(clk), .rst(rst), .q(c475ibus), .r(c475obus));
wire [temp_w*6-1:0] c476ibus;
wire [data_w*6-1:0] c476obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU476 ( .en(en), .clk(clk), .rst(rst), .q(c476ibus), .r(c476obus));
wire [temp_w*6-1:0] c477ibus;
wire [data_w*6-1:0] c477obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU477 ( .en(en), .clk(clk), .rst(rst), .q(c477ibus), .r(c477obus));
wire [temp_w*6-1:0] c478ibus;
wire [data_w*6-1:0] c478obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU478 ( .en(en), .clk(clk), .rst(rst), .q(c478ibus), .r(c478obus));
wire [temp_w*6-1:0] c479ibus;
wire [data_w*6-1:0] c479obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU479 ( .en(en), .clk(clk), .rst(rst), .q(c479ibus), .r(c479obus));
wire [temp_w*7-1:0] c480ibus;
wire [data_w*7-1:0] c480obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU480 ( .en(en), .clk(clk), .rst(rst), .q(c480ibus), .r(c480obus));
wire [temp_w*7-1:0] c481ibus;
wire [data_w*7-1:0] c481obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU481 ( .en(en), .clk(clk), .rst(rst), .q(c481ibus), .r(c481obus));
wire [temp_w*7-1:0] c482ibus;
wire [data_w*7-1:0] c482obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU482 ( .en(en), .clk(clk), .rst(rst), .q(c482ibus), .r(c482obus));
wire [temp_w*7-1:0] c483ibus;
wire [data_w*7-1:0] c483obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU483 ( .en(en), .clk(clk), .rst(rst), .q(c483ibus), .r(c483obus));
wire [temp_w*7-1:0] c484ibus;
wire [data_w*7-1:0] c484obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU484 ( .en(en), .clk(clk), .rst(rst), .q(c484ibus), .r(c484obus));
wire [temp_w*7-1:0] c485ibus;
wire [data_w*7-1:0] c485obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU485 ( .en(en), .clk(clk), .rst(rst), .q(c485ibus), .r(c485obus));
wire [temp_w*7-1:0] c486ibus;
wire [data_w*7-1:0] c486obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU486 ( .en(en), .clk(clk), .rst(rst), .q(c486ibus), .r(c486obus));
wire [temp_w*7-1:0] c487ibus;
wire [data_w*7-1:0] c487obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU487 ( .en(en), .clk(clk), .rst(rst), .q(c487ibus), .r(c487obus));
wire [temp_w*7-1:0] c488ibus;
wire [data_w*7-1:0] c488obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU488 ( .en(en), .clk(clk), .rst(rst), .q(c488ibus), .r(c488obus));
wire [temp_w*7-1:0] c489ibus;
wire [data_w*7-1:0] c489obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU489 ( .en(en), .clk(clk), .rst(rst), .q(c489ibus), .r(c489obus));
wire [temp_w*7-1:0] c490ibus;
wire [data_w*7-1:0] c490obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU490 ( .en(en), .clk(clk), .rst(rst), .q(c490ibus), .r(c490obus));
wire [temp_w*7-1:0] c491ibus;
wire [data_w*7-1:0] c491obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU491 ( .en(en), .clk(clk), .rst(rst), .q(c491ibus), .r(c491obus));
wire [temp_w*7-1:0] c492ibus;
wire [data_w*7-1:0] c492obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU492 ( .en(en), .clk(clk), .rst(rst), .q(c492ibus), .r(c492obus));
wire [temp_w*7-1:0] c493ibus;
wire [data_w*7-1:0] c493obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU493 ( .en(en), .clk(clk), .rst(rst), .q(c493ibus), .r(c493obus));
wire [temp_w*7-1:0] c494ibus;
wire [data_w*7-1:0] c494obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU494 ( .en(en), .clk(clk), .rst(rst), .q(c494ibus), .r(c494obus));
wire [temp_w*7-1:0] c495ibus;
wire [data_w*7-1:0] c495obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU495 ( .en(en), .clk(clk), .rst(rst), .q(c495ibus), .r(c495obus));
wire [temp_w*7-1:0] c496ibus;
wire [data_w*7-1:0] c496obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU496 ( .en(en), .clk(clk), .rst(rst), .q(c496ibus), .r(c496obus));
wire [temp_w*7-1:0] c497ibus;
wire [data_w*7-1:0] c497obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU497 ( .en(en), .clk(clk), .rst(rst), .q(c497ibus), .r(c497obus));
wire [temp_w*7-1:0] c498ibus;
wire [data_w*7-1:0] c498obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU498 ( .en(en), .clk(clk), .rst(rst), .q(c498ibus), .r(c498obus));
wire [temp_w*7-1:0] c499ibus;
wire [data_w*7-1:0] c499obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU499 ( .en(en), .clk(clk), .rst(rst), .q(c499ibus), .r(c499obus));
wire [temp_w*7-1:0] c500ibus;
wire [data_w*7-1:0] c500obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU500 ( .en(en), .clk(clk), .rst(rst), .q(c500ibus), .r(c500obus));
wire [temp_w*7-1:0] c501ibus;
wire [data_w*7-1:0] c501obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU501 ( .en(en), .clk(clk), .rst(rst), .q(c501ibus), .r(c501obus));
wire [temp_w*7-1:0] c502ibus;
wire [data_w*7-1:0] c502obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU502 ( .en(en), .clk(clk), .rst(rst), .q(c502ibus), .r(c502obus));
wire [temp_w*7-1:0] c503ibus;
wire [data_w*7-1:0] c503obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU503 ( .en(en), .clk(clk), .rst(rst), .q(c503ibus), .r(c503obus));
wire [temp_w*7-1:0] c504ibus;
wire [data_w*7-1:0] c504obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU504 ( .en(en), .clk(clk), .rst(rst), .q(c504ibus), .r(c504obus));
wire [temp_w*7-1:0] c505ibus;
wire [data_w*7-1:0] c505obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU505 ( .en(en), .clk(clk), .rst(rst), .q(c505ibus), .r(c505obus));
wire [temp_w*7-1:0] c506ibus;
wire [data_w*7-1:0] c506obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU506 ( .en(en), .clk(clk), .rst(rst), .q(c506ibus), .r(c506obus));
wire [temp_w*7-1:0] c507ibus;
wire [data_w*7-1:0] c507obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU507 ( .en(en), .clk(clk), .rst(rst), .q(c507ibus), .r(c507obus));
wire [temp_w*7-1:0] c508ibus;
wire [data_w*7-1:0] c508obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU508 ( .en(en), .clk(clk), .rst(rst), .q(c508ibus), .r(c508obus));
wire [temp_w*7-1:0] c509ibus;
wire [data_w*7-1:0] c509obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU509 ( .en(en), .clk(clk), .rst(rst), .q(c509ibus), .r(c509obus));
wire [temp_w*7-1:0] c510ibus;
wire [data_w*7-1:0] c510obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU510 ( .en(en), .clk(clk), .rst(rst), .q(c510ibus), .r(c510obus));
wire [temp_w*7-1:0] c511ibus;
wire [data_w*7-1:0] c511obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU511 ( .en(en), .clk(clk), .rst(rst), .q(c511ibus), .r(c511obus));
wire [temp_w*7-1:0] c512ibus;
wire [data_w*7-1:0] c512obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU512 ( .en(en), .clk(clk), .rst(rst), .q(c512ibus), .r(c512obus));
wire [temp_w*7-1:0] c513ibus;
wire [data_w*7-1:0] c513obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU513 ( .en(en), .clk(clk), .rst(rst), .q(c513ibus), .r(c513obus));
wire [temp_w*7-1:0] c514ibus;
wire [data_w*7-1:0] c514obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU514 ( .en(en), .clk(clk), .rst(rst), .q(c514ibus), .r(c514obus));
wire [temp_w*7-1:0] c515ibus;
wire [data_w*7-1:0] c515obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU515 ( .en(en), .clk(clk), .rst(rst), .q(c515ibus), .r(c515obus));
wire [temp_w*7-1:0] c516ibus;
wire [data_w*7-1:0] c516obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU516 ( .en(en), .clk(clk), .rst(rst), .q(c516ibus), .r(c516obus));
wire [temp_w*7-1:0] c517ibus;
wire [data_w*7-1:0] c517obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU517 ( .en(en), .clk(clk), .rst(rst), .q(c517ibus), .r(c517obus));
wire [temp_w*7-1:0] c518ibus;
wire [data_w*7-1:0] c518obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU518 ( .en(en), .clk(clk), .rst(rst), .q(c518ibus), .r(c518obus));
wire [temp_w*7-1:0] c519ibus;
wire [data_w*7-1:0] c519obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU519 ( .en(en), .clk(clk), .rst(rst), .q(c519ibus), .r(c519obus));
wire [temp_w*7-1:0] c520ibus;
wire [data_w*7-1:0] c520obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU520 ( .en(en), .clk(clk), .rst(rst), .q(c520ibus), .r(c520obus));
wire [temp_w*7-1:0] c521ibus;
wire [data_w*7-1:0] c521obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU521 ( .en(en), .clk(clk), .rst(rst), .q(c521ibus), .r(c521obus));
wire [temp_w*7-1:0] c522ibus;
wire [data_w*7-1:0] c522obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU522 ( .en(en), .clk(clk), .rst(rst), .q(c522ibus), .r(c522obus));
wire [temp_w*7-1:0] c523ibus;
wire [data_w*7-1:0] c523obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU523 ( .en(en), .clk(clk), .rst(rst), .q(c523ibus), .r(c523obus));
wire [temp_w*7-1:0] c524ibus;
wire [data_w*7-1:0] c524obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU524 ( .en(en), .clk(clk), .rst(rst), .q(c524ibus), .r(c524obus));
wire [temp_w*7-1:0] c525ibus;
wire [data_w*7-1:0] c525obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU525 ( .en(en), .clk(clk), .rst(rst), .q(c525ibus), .r(c525obus));
wire [temp_w*7-1:0] c526ibus;
wire [data_w*7-1:0] c526obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU526 ( .en(en), .clk(clk), .rst(rst), .q(c526ibus), .r(c526obus));
wire [temp_w*7-1:0] c527ibus;
wire [data_w*7-1:0] c527obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU527 ( .en(en), .clk(clk), .rst(rst), .q(c527ibus), .r(c527obus));
wire [temp_w*7-1:0] c528ibus;
wire [data_w*7-1:0] c528obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU528 ( .en(en), .clk(clk), .rst(rst), .q(c528ibus), .r(c528obus));
wire [temp_w*7-1:0] c529ibus;
wire [data_w*7-1:0] c529obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU529 ( .en(en), .clk(clk), .rst(rst), .q(c529ibus), .r(c529obus));
wire [temp_w*7-1:0] c530ibus;
wire [data_w*7-1:0] c530obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU530 ( .en(en), .clk(clk), .rst(rst), .q(c530ibus), .r(c530obus));
wire [temp_w*7-1:0] c531ibus;
wire [data_w*7-1:0] c531obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU531 ( .en(en), .clk(clk), .rst(rst), .q(c531ibus), .r(c531obus));
wire [temp_w*7-1:0] c532ibus;
wire [data_w*7-1:0] c532obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU532 ( .en(en), .clk(clk), .rst(rst), .q(c532ibus), .r(c532obus));
wire [temp_w*7-1:0] c533ibus;
wire [data_w*7-1:0] c533obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU533 ( .en(en), .clk(clk), .rst(rst), .q(c533ibus), .r(c533obus));
wire [temp_w*7-1:0] c534ibus;
wire [data_w*7-1:0] c534obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU534 ( .en(en), .clk(clk), .rst(rst), .q(c534ibus), .r(c534obus));
wire [temp_w*7-1:0] c535ibus;
wire [data_w*7-1:0] c535obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU535 ( .en(en), .clk(clk), .rst(rst), .q(c535ibus), .r(c535obus));
wire [temp_w*7-1:0] c536ibus;
wire [data_w*7-1:0] c536obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU536 ( .en(en), .clk(clk), .rst(rst), .q(c536ibus), .r(c536obus));
wire [temp_w*7-1:0] c537ibus;
wire [data_w*7-1:0] c537obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU537 ( .en(en), .clk(clk), .rst(rst), .q(c537ibus), .r(c537obus));
wire [temp_w*7-1:0] c538ibus;
wire [data_w*7-1:0] c538obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU538 ( .en(en), .clk(clk), .rst(rst), .q(c538ibus), .r(c538obus));
wire [temp_w*7-1:0] c539ibus;
wire [data_w*7-1:0] c539obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU539 ( .en(en), .clk(clk), .rst(rst), .q(c539ibus), .r(c539obus));
wire [temp_w*7-1:0] c540ibus;
wire [data_w*7-1:0] c540obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU540 ( .en(en), .clk(clk), .rst(rst), .q(c540ibus), .r(c540obus));
wire [temp_w*7-1:0] c541ibus;
wire [data_w*7-1:0] c541obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU541 ( .en(en), .clk(clk), .rst(rst), .q(c541ibus), .r(c541obus));
wire [temp_w*7-1:0] c542ibus;
wire [data_w*7-1:0] c542obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU542 ( .en(en), .clk(clk), .rst(rst), .q(c542ibus), .r(c542obus));
wire [temp_w*7-1:0] c543ibus;
wire [data_w*7-1:0] c543obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU543 ( .en(en), .clk(clk), .rst(rst), .q(c543ibus), .r(c543obus));
wire [temp_w*7-1:0] c544ibus;
wire [data_w*7-1:0] c544obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU544 ( .en(en), .clk(clk), .rst(rst), .q(c544ibus), .r(c544obus));
wire [temp_w*7-1:0] c545ibus;
wire [data_w*7-1:0] c545obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU545 ( .en(en), .clk(clk), .rst(rst), .q(c545ibus), .r(c545obus));
wire [temp_w*7-1:0] c546ibus;
wire [data_w*7-1:0] c546obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU546 ( .en(en), .clk(clk), .rst(rst), .q(c546ibus), .r(c546obus));
wire [temp_w*7-1:0] c547ibus;
wire [data_w*7-1:0] c547obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU547 ( .en(en), .clk(clk), .rst(rst), .q(c547ibus), .r(c547obus));
wire [temp_w*7-1:0] c548ibus;
wire [data_w*7-1:0] c548obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU548 ( .en(en), .clk(clk), .rst(rst), .q(c548ibus), .r(c548obus));
wire [temp_w*7-1:0] c549ibus;
wire [data_w*7-1:0] c549obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU549 ( .en(en), .clk(clk), .rst(rst), .q(c549ibus), .r(c549obus));
wire [temp_w*7-1:0] c550ibus;
wire [data_w*7-1:0] c550obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU550 ( .en(en), .clk(clk), .rst(rst), .q(c550ibus), .r(c550obus));
wire [temp_w*7-1:0] c551ibus;
wire [data_w*7-1:0] c551obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU551 ( .en(en), .clk(clk), .rst(rst), .q(c551ibus), .r(c551obus));
wire [temp_w*7-1:0] c552ibus;
wire [data_w*7-1:0] c552obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU552 ( .en(en), .clk(clk), .rst(rst), .q(c552ibus), .r(c552obus));
wire [temp_w*7-1:0] c553ibus;
wire [data_w*7-1:0] c553obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU553 ( .en(en), .clk(clk), .rst(rst), .q(c553ibus), .r(c553obus));
wire [temp_w*7-1:0] c554ibus;
wire [data_w*7-1:0] c554obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU554 ( .en(en), .clk(clk), .rst(rst), .q(c554ibus), .r(c554obus));
wire [temp_w*7-1:0] c555ibus;
wire [data_w*7-1:0] c555obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU555 ( .en(en), .clk(clk), .rst(rst), .q(c555ibus), .r(c555obus));
wire [temp_w*7-1:0] c556ibus;
wire [data_w*7-1:0] c556obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU556 ( .en(en), .clk(clk), .rst(rst), .q(c556ibus), .r(c556obus));
wire [temp_w*7-1:0] c557ibus;
wire [data_w*7-1:0] c557obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU557 ( .en(en), .clk(clk), .rst(rst), .q(c557ibus), .r(c557obus));
wire [temp_w*7-1:0] c558ibus;
wire [data_w*7-1:0] c558obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU558 ( .en(en), .clk(clk), .rst(rst), .q(c558ibus), .r(c558obus));
wire [temp_w*7-1:0] c559ibus;
wire [data_w*7-1:0] c559obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU559 ( .en(en), .clk(clk), .rst(rst), .q(c559ibus), .r(c559obus));
wire [temp_w*7-1:0] c560ibus;
wire [data_w*7-1:0] c560obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU560 ( .en(en), .clk(clk), .rst(rst), .q(c560ibus), .r(c560obus));
wire [temp_w*7-1:0] c561ibus;
wire [data_w*7-1:0] c561obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU561 ( .en(en), .clk(clk), .rst(rst), .q(c561ibus), .r(c561obus));
wire [temp_w*7-1:0] c562ibus;
wire [data_w*7-1:0] c562obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU562 ( .en(en), .clk(clk), .rst(rst), .q(c562ibus), .r(c562obus));
wire [temp_w*7-1:0] c563ibus;
wire [data_w*7-1:0] c563obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU563 ( .en(en), .clk(clk), .rst(rst), .q(c563ibus), .r(c563obus));
wire [temp_w*7-1:0] c564ibus;
wire [data_w*7-1:0] c564obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU564 ( .en(en), .clk(clk), .rst(rst), .q(c564ibus), .r(c564obus));
wire [temp_w*7-1:0] c565ibus;
wire [data_w*7-1:0] c565obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU565 ( .en(en), .clk(clk), .rst(rst), .q(c565ibus), .r(c565obus));
wire [temp_w*7-1:0] c566ibus;
wire [data_w*7-1:0] c566obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU566 ( .en(en), .clk(clk), .rst(rst), .q(c566ibus), .r(c566obus));
wire [temp_w*7-1:0] c567ibus;
wire [data_w*7-1:0] c567obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU567 ( .en(en), .clk(clk), .rst(rst), .q(c567ibus), .r(c567obus));
wire [temp_w*7-1:0] c568ibus;
wire [data_w*7-1:0] c568obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU568 ( .en(en), .clk(clk), .rst(rst), .q(c568ibus), .r(c568obus));
wire [temp_w*7-1:0] c569ibus;
wire [data_w*7-1:0] c569obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU569 ( .en(en), .clk(clk), .rst(rst), .q(c569ibus), .r(c569obus));
wire [temp_w*7-1:0] c570ibus;
wire [data_w*7-1:0] c570obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU570 ( .en(en), .clk(clk), .rst(rst), .q(c570ibus), .r(c570obus));
wire [temp_w*7-1:0] c571ibus;
wire [data_w*7-1:0] c571obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU571 ( .en(en), .clk(clk), .rst(rst), .q(c571ibus), .r(c571obus));
wire [temp_w*7-1:0] c572ibus;
wire [data_w*7-1:0] c572obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU572 ( .en(en), .clk(clk), .rst(rst), .q(c572ibus), .r(c572obus));
wire [temp_w*7-1:0] c573ibus;
wire [data_w*7-1:0] c573obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU573 ( .en(en), .clk(clk), .rst(rst), .q(c573ibus), .r(c573obus));
wire [temp_w*7-1:0] c574ibus;
wire [data_w*7-1:0] c574obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU574 ( .en(en), .clk(clk), .rst(rst), .q(c574ibus), .r(c574obus));
wire [temp_w*7-1:0] c575ibus;
wire [data_w*7-1:0] c575obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU575 ( .en(en), .clk(clk), .rst(rst), .q(c575ibus), .r(c575obus));
wire [temp_w*6-1:0] c576ibus;
wire [data_w*6-1:0] c576obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU576 ( .en(en), .clk(clk), .rst(rst), .q(c576ibus), .r(c576obus));
wire [temp_w*6-1:0] c577ibus;
wire [data_w*6-1:0] c577obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU577 ( .en(en), .clk(clk), .rst(rst), .q(c577ibus), .r(c577obus));
wire [temp_w*6-1:0] c578ibus;
wire [data_w*6-1:0] c578obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU578 ( .en(en), .clk(clk), .rst(rst), .q(c578ibus), .r(c578obus));
wire [temp_w*6-1:0] c579ibus;
wire [data_w*6-1:0] c579obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU579 ( .en(en), .clk(clk), .rst(rst), .q(c579ibus), .r(c579obus));
wire [temp_w*6-1:0] c580ibus;
wire [data_w*6-1:0] c580obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU580 ( .en(en), .clk(clk), .rst(rst), .q(c580ibus), .r(c580obus));
wire [temp_w*6-1:0] c581ibus;
wire [data_w*6-1:0] c581obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU581 ( .en(en), .clk(clk), .rst(rst), .q(c581ibus), .r(c581obus));
wire [temp_w*6-1:0] c582ibus;
wire [data_w*6-1:0] c582obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU582 ( .en(en), .clk(clk), .rst(rst), .q(c582ibus), .r(c582obus));
wire [temp_w*6-1:0] c583ibus;
wire [data_w*6-1:0] c583obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU583 ( .en(en), .clk(clk), .rst(rst), .q(c583ibus), .r(c583obus));
wire [temp_w*6-1:0] c584ibus;
wire [data_w*6-1:0] c584obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU584 ( .en(en), .clk(clk), .rst(rst), .q(c584ibus), .r(c584obus));
wire [temp_w*6-1:0] c585ibus;
wire [data_w*6-1:0] c585obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU585 ( .en(en), .clk(clk), .rst(rst), .q(c585ibus), .r(c585obus));
wire [temp_w*6-1:0] c586ibus;
wire [data_w*6-1:0] c586obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU586 ( .en(en), .clk(clk), .rst(rst), .q(c586ibus), .r(c586obus));
wire [temp_w*6-1:0] c587ibus;
wire [data_w*6-1:0] c587obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU587 ( .en(en), .clk(clk), .rst(rst), .q(c587ibus), .r(c587obus));
wire [temp_w*6-1:0] c588ibus;
wire [data_w*6-1:0] c588obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU588 ( .en(en), .clk(clk), .rst(rst), .q(c588ibus), .r(c588obus));
wire [temp_w*6-1:0] c589ibus;
wire [data_w*6-1:0] c589obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU589 ( .en(en), .clk(clk), .rst(rst), .q(c589ibus), .r(c589obus));
wire [temp_w*6-1:0] c590ibus;
wire [data_w*6-1:0] c590obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU590 ( .en(en), .clk(clk), .rst(rst), .q(c590ibus), .r(c590obus));
wire [temp_w*6-1:0] c591ibus;
wire [data_w*6-1:0] c591obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU591 ( .en(en), .clk(clk), .rst(rst), .q(c591ibus), .r(c591obus));
wire [temp_w*6-1:0] c592ibus;
wire [data_w*6-1:0] c592obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU592 ( .en(en), .clk(clk), .rst(rst), .q(c592ibus), .r(c592obus));
wire [temp_w*6-1:0] c593ibus;
wire [data_w*6-1:0] c593obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU593 ( .en(en), .clk(clk), .rst(rst), .q(c593ibus), .r(c593obus));
wire [temp_w*6-1:0] c594ibus;
wire [data_w*6-1:0] c594obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU594 ( .en(en), .clk(clk), .rst(rst), .q(c594ibus), .r(c594obus));
wire [temp_w*6-1:0] c595ibus;
wire [data_w*6-1:0] c595obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU595 ( .en(en), .clk(clk), .rst(rst), .q(c595ibus), .r(c595obus));
wire [temp_w*6-1:0] c596ibus;
wire [data_w*6-1:0] c596obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU596 ( .en(en), .clk(clk), .rst(rst), .q(c596ibus), .r(c596obus));
wire [temp_w*6-1:0] c597ibus;
wire [data_w*6-1:0] c597obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU597 ( .en(en), .clk(clk), .rst(rst), .q(c597ibus), .r(c597obus));
wire [temp_w*6-1:0] c598ibus;
wire [data_w*6-1:0] c598obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU598 ( .en(en), .clk(clk), .rst(rst), .q(c598ibus), .r(c598obus));
wire [temp_w*6-1:0] c599ibus;
wire [data_w*6-1:0] c599obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU599 ( .en(en), .clk(clk), .rst(rst), .q(c599ibus), .r(c599obus));
wire [temp_w*6-1:0] c600ibus;
wire [data_w*6-1:0] c600obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU600 ( .en(en), .clk(clk), .rst(rst), .q(c600ibus), .r(c600obus));
wire [temp_w*6-1:0] c601ibus;
wire [data_w*6-1:0] c601obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU601 ( .en(en), .clk(clk), .rst(rst), .q(c601ibus), .r(c601obus));
wire [temp_w*6-1:0] c602ibus;
wire [data_w*6-1:0] c602obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU602 ( .en(en), .clk(clk), .rst(rst), .q(c602ibus), .r(c602obus));
wire [temp_w*6-1:0] c603ibus;
wire [data_w*6-1:0] c603obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU603 ( .en(en), .clk(clk), .rst(rst), .q(c603ibus), .r(c603obus));
wire [temp_w*6-1:0] c604ibus;
wire [data_w*6-1:0] c604obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU604 ( .en(en), .clk(clk), .rst(rst), .q(c604ibus), .r(c604obus));
wire [temp_w*6-1:0] c605ibus;
wire [data_w*6-1:0] c605obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU605 ( .en(en), .clk(clk), .rst(rst), .q(c605ibus), .r(c605obus));
wire [temp_w*6-1:0] c606ibus;
wire [data_w*6-1:0] c606obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU606 ( .en(en), .clk(clk), .rst(rst), .q(c606ibus), .r(c606obus));
wire [temp_w*6-1:0] c607ibus;
wire [data_w*6-1:0] c607obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU607 ( .en(en), .clk(clk), .rst(rst), .q(c607ibus), .r(c607obus));
wire [temp_w*6-1:0] c608ibus;
wire [data_w*6-1:0] c608obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU608 ( .en(en), .clk(clk), .rst(rst), .q(c608ibus), .r(c608obus));
wire [temp_w*6-1:0] c609ibus;
wire [data_w*6-1:0] c609obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU609 ( .en(en), .clk(clk), .rst(rst), .q(c609ibus), .r(c609obus));
wire [temp_w*6-1:0] c610ibus;
wire [data_w*6-1:0] c610obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU610 ( .en(en), .clk(clk), .rst(rst), .q(c610ibus), .r(c610obus));
wire [temp_w*6-1:0] c611ibus;
wire [data_w*6-1:0] c611obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU611 ( .en(en), .clk(clk), .rst(rst), .q(c611ibus), .r(c611obus));
wire [temp_w*6-1:0] c612ibus;
wire [data_w*6-1:0] c612obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU612 ( .en(en), .clk(clk), .rst(rst), .q(c612ibus), .r(c612obus));
wire [temp_w*6-1:0] c613ibus;
wire [data_w*6-1:0] c613obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU613 ( .en(en), .clk(clk), .rst(rst), .q(c613ibus), .r(c613obus));
wire [temp_w*6-1:0] c614ibus;
wire [data_w*6-1:0] c614obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU614 ( .en(en), .clk(clk), .rst(rst), .q(c614ibus), .r(c614obus));
wire [temp_w*6-1:0] c615ibus;
wire [data_w*6-1:0] c615obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU615 ( .en(en), .clk(clk), .rst(rst), .q(c615ibus), .r(c615obus));
wire [temp_w*6-1:0] c616ibus;
wire [data_w*6-1:0] c616obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU616 ( .en(en), .clk(clk), .rst(rst), .q(c616ibus), .r(c616obus));
wire [temp_w*6-1:0] c617ibus;
wire [data_w*6-1:0] c617obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU617 ( .en(en), .clk(clk), .rst(rst), .q(c617ibus), .r(c617obus));
wire [temp_w*6-1:0] c618ibus;
wire [data_w*6-1:0] c618obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU618 ( .en(en), .clk(clk), .rst(rst), .q(c618ibus), .r(c618obus));
wire [temp_w*6-1:0] c619ibus;
wire [data_w*6-1:0] c619obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU619 ( .en(en), .clk(clk), .rst(rst), .q(c619ibus), .r(c619obus));
wire [temp_w*6-1:0] c620ibus;
wire [data_w*6-1:0] c620obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU620 ( .en(en), .clk(clk), .rst(rst), .q(c620ibus), .r(c620obus));
wire [temp_w*6-1:0] c621ibus;
wire [data_w*6-1:0] c621obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU621 ( .en(en), .clk(clk), .rst(rst), .q(c621ibus), .r(c621obus));
wire [temp_w*6-1:0] c622ibus;
wire [data_w*6-1:0] c622obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU622 ( .en(en), .clk(clk), .rst(rst), .q(c622ibus), .r(c622obus));
wire [temp_w*6-1:0] c623ibus;
wire [data_w*6-1:0] c623obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU623 ( .en(en), .clk(clk), .rst(rst), .q(c623ibus), .r(c623obus));
wire [temp_w*6-1:0] c624ibus;
wire [data_w*6-1:0] c624obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU624 ( .en(en), .clk(clk), .rst(rst), .q(c624ibus), .r(c624obus));
wire [temp_w*6-1:0] c625ibus;
wire [data_w*6-1:0] c625obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU625 ( .en(en), .clk(clk), .rst(rst), .q(c625ibus), .r(c625obus));
wire [temp_w*6-1:0] c626ibus;
wire [data_w*6-1:0] c626obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU626 ( .en(en), .clk(clk), .rst(rst), .q(c626ibus), .r(c626obus));
wire [temp_w*6-1:0] c627ibus;
wire [data_w*6-1:0] c627obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU627 ( .en(en), .clk(clk), .rst(rst), .q(c627ibus), .r(c627obus));
wire [temp_w*6-1:0] c628ibus;
wire [data_w*6-1:0] c628obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU628 ( .en(en), .clk(clk), .rst(rst), .q(c628ibus), .r(c628obus));
wire [temp_w*6-1:0] c629ibus;
wire [data_w*6-1:0] c629obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU629 ( .en(en), .clk(clk), .rst(rst), .q(c629ibus), .r(c629obus));
wire [temp_w*6-1:0] c630ibus;
wire [data_w*6-1:0] c630obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU630 ( .en(en), .clk(clk), .rst(rst), .q(c630ibus), .r(c630obus));
wire [temp_w*6-1:0] c631ibus;
wire [data_w*6-1:0] c631obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU631 ( .en(en), .clk(clk), .rst(rst), .q(c631ibus), .r(c631obus));
wire [temp_w*6-1:0] c632ibus;
wire [data_w*6-1:0] c632obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU632 ( .en(en), .clk(clk), .rst(rst), .q(c632ibus), .r(c632obus));
wire [temp_w*6-1:0] c633ibus;
wire [data_w*6-1:0] c633obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU633 ( .en(en), .clk(clk), .rst(rst), .q(c633ibus), .r(c633obus));
wire [temp_w*6-1:0] c634ibus;
wire [data_w*6-1:0] c634obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU634 ( .en(en), .clk(clk), .rst(rst), .q(c634ibus), .r(c634obus));
wire [temp_w*6-1:0] c635ibus;
wire [data_w*6-1:0] c635obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU635 ( .en(en), .clk(clk), .rst(rst), .q(c635ibus), .r(c635obus));
wire [temp_w*6-1:0] c636ibus;
wire [data_w*6-1:0] c636obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU636 ( .en(en), .clk(clk), .rst(rst), .q(c636ibus), .r(c636obus));
wire [temp_w*6-1:0] c637ibus;
wire [data_w*6-1:0] c637obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU637 ( .en(en), .clk(clk), .rst(rst), .q(c637ibus), .r(c637obus));
wire [temp_w*6-1:0] c638ibus;
wire [data_w*6-1:0] c638obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU638 ( .en(en), .clk(clk), .rst(rst), .q(c638ibus), .r(c638obus));
wire [temp_w*6-1:0] c639ibus;
wire [data_w*6-1:0] c639obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU639 ( .en(en), .clk(clk), .rst(rst), .q(c639ibus), .r(c639obus));
wire [temp_w*6-1:0] c640ibus;
wire [data_w*6-1:0] c640obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU640 ( .en(en), .clk(clk), .rst(rst), .q(c640ibus), .r(c640obus));
wire [temp_w*6-1:0] c641ibus;
wire [data_w*6-1:0] c641obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU641 ( .en(en), .clk(clk), .rst(rst), .q(c641ibus), .r(c641obus));
wire [temp_w*6-1:0] c642ibus;
wire [data_w*6-1:0] c642obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU642 ( .en(en), .clk(clk), .rst(rst), .q(c642ibus), .r(c642obus));
wire [temp_w*6-1:0] c643ibus;
wire [data_w*6-1:0] c643obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU643 ( .en(en), .clk(clk), .rst(rst), .q(c643ibus), .r(c643obus));
wire [temp_w*6-1:0] c644ibus;
wire [data_w*6-1:0] c644obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU644 ( .en(en), .clk(clk), .rst(rst), .q(c644ibus), .r(c644obus));
wire [temp_w*6-1:0] c645ibus;
wire [data_w*6-1:0] c645obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU645 ( .en(en), .clk(clk), .rst(rst), .q(c645ibus), .r(c645obus));
wire [temp_w*6-1:0] c646ibus;
wire [data_w*6-1:0] c646obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU646 ( .en(en), .clk(clk), .rst(rst), .q(c646ibus), .r(c646obus));
wire [temp_w*6-1:0] c647ibus;
wire [data_w*6-1:0] c647obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU647 ( .en(en), .clk(clk), .rst(rst), .q(c647ibus), .r(c647obus));
wire [temp_w*6-1:0] c648ibus;
wire [data_w*6-1:0] c648obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU648 ( .en(en), .clk(clk), .rst(rst), .q(c648ibus), .r(c648obus));
wire [temp_w*6-1:0] c649ibus;
wire [data_w*6-1:0] c649obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU649 ( .en(en), .clk(clk), .rst(rst), .q(c649ibus), .r(c649obus));
wire [temp_w*6-1:0] c650ibus;
wire [data_w*6-1:0] c650obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU650 ( .en(en), .clk(clk), .rst(rst), .q(c650ibus), .r(c650obus));
wire [temp_w*6-1:0] c651ibus;
wire [data_w*6-1:0] c651obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU651 ( .en(en), .clk(clk), .rst(rst), .q(c651ibus), .r(c651obus));
wire [temp_w*6-1:0] c652ibus;
wire [data_w*6-1:0] c652obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU652 ( .en(en), .clk(clk), .rst(rst), .q(c652ibus), .r(c652obus));
wire [temp_w*6-1:0] c653ibus;
wire [data_w*6-1:0] c653obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU653 ( .en(en), .clk(clk), .rst(rst), .q(c653ibus), .r(c653obus));
wire [temp_w*6-1:0] c654ibus;
wire [data_w*6-1:0] c654obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU654 ( .en(en), .clk(clk), .rst(rst), .q(c654ibus), .r(c654obus));
wire [temp_w*6-1:0] c655ibus;
wire [data_w*6-1:0] c655obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU655 ( .en(en), .clk(clk), .rst(rst), .q(c655ibus), .r(c655obus));
wire [temp_w*6-1:0] c656ibus;
wire [data_w*6-1:0] c656obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU656 ( .en(en), .clk(clk), .rst(rst), .q(c656ibus), .r(c656obus));
wire [temp_w*6-1:0] c657ibus;
wire [data_w*6-1:0] c657obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU657 ( .en(en), .clk(clk), .rst(rst), .q(c657ibus), .r(c657obus));
wire [temp_w*6-1:0] c658ibus;
wire [data_w*6-1:0] c658obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU658 ( .en(en), .clk(clk), .rst(rst), .q(c658ibus), .r(c658obus));
wire [temp_w*6-1:0] c659ibus;
wire [data_w*6-1:0] c659obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU659 ( .en(en), .clk(clk), .rst(rst), .q(c659ibus), .r(c659obus));
wire [temp_w*6-1:0] c660ibus;
wire [data_w*6-1:0] c660obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU660 ( .en(en), .clk(clk), .rst(rst), .q(c660ibus), .r(c660obus));
wire [temp_w*6-1:0] c661ibus;
wire [data_w*6-1:0] c661obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU661 ( .en(en), .clk(clk), .rst(rst), .q(c661ibus), .r(c661obus));
wire [temp_w*6-1:0] c662ibus;
wire [data_w*6-1:0] c662obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU662 ( .en(en), .clk(clk), .rst(rst), .q(c662ibus), .r(c662obus));
wire [temp_w*6-1:0] c663ibus;
wire [data_w*6-1:0] c663obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU663 ( .en(en), .clk(clk), .rst(rst), .q(c663ibus), .r(c663obus));
wire [temp_w*6-1:0] c664ibus;
wire [data_w*6-1:0] c664obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU664 ( .en(en), .clk(clk), .rst(rst), .q(c664ibus), .r(c664obus));
wire [temp_w*6-1:0] c665ibus;
wire [data_w*6-1:0] c665obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU665 ( .en(en), .clk(clk), .rst(rst), .q(c665ibus), .r(c665obus));
wire [temp_w*6-1:0] c666ibus;
wire [data_w*6-1:0] c666obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU666 ( .en(en), .clk(clk), .rst(rst), .q(c666ibus), .r(c666obus));
wire [temp_w*6-1:0] c667ibus;
wire [data_w*6-1:0] c667obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU667 ( .en(en), .clk(clk), .rst(rst), .q(c667ibus), .r(c667obus));
wire [temp_w*6-1:0] c668ibus;
wire [data_w*6-1:0] c668obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU668 ( .en(en), .clk(clk), .rst(rst), .q(c668ibus), .r(c668obus));
wire [temp_w*6-1:0] c669ibus;
wire [data_w*6-1:0] c669obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU669 ( .en(en), .clk(clk), .rst(rst), .q(c669ibus), .r(c669obus));
wire [temp_w*6-1:0] c670ibus;
wire [data_w*6-1:0] c670obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU670 ( .en(en), .clk(clk), .rst(rst), .q(c670ibus), .r(c670obus));
wire [temp_w*6-1:0] c671ibus;
wire [data_w*6-1:0] c671obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU671 ( .en(en), .clk(clk), .rst(rst), .q(c671ibus), .r(c671obus));
wire [temp_w*6-1:0] c672ibus;
wire [data_w*6-1:0] c672obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU672 ( .en(en), .clk(clk), .rst(rst), .q(c672ibus), .r(c672obus));
wire [temp_w*6-1:0] c673ibus;
wire [data_w*6-1:0] c673obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU673 ( .en(en), .clk(clk), .rst(rst), .q(c673ibus), .r(c673obus));
wire [temp_w*6-1:0] c674ibus;
wire [data_w*6-1:0] c674obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU674 ( .en(en), .clk(clk), .rst(rst), .q(c674ibus), .r(c674obus));
wire [temp_w*6-1:0] c675ibus;
wire [data_w*6-1:0] c675obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU675 ( .en(en), .clk(clk), .rst(rst), .q(c675ibus), .r(c675obus));
wire [temp_w*6-1:0] c676ibus;
wire [data_w*6-1:0] c676obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU676 ( .en(en), .clk(clk), .rst(rst), .q(c676ibus), .r(c676obus));
wire [temp_w*6-1:0] c677ibus;
wire [data_w*6-1:0] c677obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU677 ( .en(en), .clk(clk), .rst(rst), .q(c677ibus), .r(c677obus));
wire [temp_w*6-1:0] c678ibus;
wire [data_w*6-1:0] c678obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU678 ( .en(en), .clk(clk), .rst(rst), .q(c678ibus), .r(c678obus));
wire [temp_w*6-1:0] c679ibus;
wire [data_w*6-1:0] c679obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU679 ( .en(en), .clk(clk), .rst(rst), .q(c679ibus), .r(c679obus));
wire [temp_w*6-1:0] c680ibus;
wire [data_w*6-1:0] c680obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU680 ( .en(en), .clk(clk), .rst(rst), .q(c680ibus), .r(c680obus));
wire [temp_w*6-1:0] c681ibus;
wire [data_w*6-1:0] c681obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU681 ( .en(en), .clk(clk), .rst(rst), .q(c681ibus), .r(c681obus));
wire [temp_w*6-1:0] c682ibus;
wire [data_w*6-1:0] c682obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU682 ( .en(en), .clk(clk), .rst(rst), .q(c682ibus), .r(c682obus));
wire [temp_w*6-1:0] c683ibus;
wire [data_w*6-1:0] c683obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU683 ( .en(en), .clk(clk), .rst(rst), .q(c683ibus), .r(c683obus));
wire [temp_w*6-1:0] c684ibus;
wire [data_w*6-1:0] c684obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU684 ( .en(en), .clk(clk), .rst(rst), .q(c684ibus), .r(c684obus));
wire [temp_w*6-1:0] c685ibus;
wire [data_w*6-1:0] c685obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU685 ( .en(en), .clk(clk), .rst(rst), .q(c685ibus), .r(c685obus));
wire [temp_w*6-1:0] c686ibus;
wire [data_w*6-1:0] c686obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU686 ( .en(en), .clk(clk), .rst(rst), .q(c686ibus), .r(c686obus));
wire [temp_w*6-1:0] c687ibus;
wire [data_w*6-1:0] c687obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU687 ( .en(en), .clk(clk), .rst(rst), .q(c687ibus), .r(c687obus));
wire [temp_w*6-1:0] c688ibus;
wire [data_w*6-1:0] c688obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU688 ( .en(en), .clk(clk), .rst(rst), .q(c688ibus), .r(c688obus));
wire [temp_w*6-1:0] c689ibus;
wire [data_w*6-1:0] c689obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU689 ( .en(en), .clk(clk), .rst(rst), .q(c689ibus), .r(c689obus));
wire [temp_w*6-1:0] c690ibus;
wire [data_w*6-1:0] c690obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU690 ( .en(en), .clk(clk), .rst(rst), .q(c690ibus), .r(c690obus));
wire [temp_w*6-1:0] c691ibus;
wire [data_w*6-1:0] c691obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU691 ( .en(en), .clk(clk), .rst(rst), .q(c691ibus), .r(c691obus));
wire [temp_w*6-1:0] c692ibus;
wire [data_w*6-1:0] c692obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU692 ( .en(en), .clk(clk), .rst(rst), .q(c692ibus), .r(c692obus));
wire [temp_w*6-1:0] c693ibus;
wire [data_w*6-1:0] c693obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU693 ( .en(en), .clk(clk), .rst(rst), .q(c693ibus), .r(c693obus));
wire [temp_w*6-1:0] c694ibus;
wire [data_w*6-1:0] c694obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU694 ( .en(en), .clk(clk), .rst(rst), .q(c694ibus), .r(c694obus));
wire [temp_w*6-1:0] c695ibus;
wire [data_w*6-1:0] c695obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU695 ( .en(en), .clk(clk), .rst(rst), .q(c695ibus), .r(c695obus));
wire [temp_w*6-1:0] c696ibus;
wire [data_w*6-1:0] c696obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU696 ( .en(en), .clk(clk), .rst(rst), .q(c696ibus), .r(c696obus));
wire [temp_w*6-1:0] c697ibus;
wire [data_w*6-1:0] c697obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU697 ( .en(en), .clk(clk), .rst(rst), .q(c697ibus), .r(c697obus));
wire [temp_w*6-1:0] c698ibus;
wire [data_w*6-1:0] c698obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU698 ( .en(en), .clk(clk), .rst(rst), .q(c698ibus), .r(c698obus));
wire [temp_w*6-1:0] c699ibus;
wire [data_w*6-1:0] c699obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU699 ( .en(en), .clk(clk), .rst(rst), .q(c699ibus), .r(c699obus));
wire [temp_w*6-1:0] c700ibus;
wire [data_w*6-1:0] c700obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU700 ( .en(en), .clk(clk), .rst(rst), .q(c700ibus), .r(c700obus));
wire [temp_w*6-1:0] c701ibus;
wire [data_w*6-1:0] c701obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU701 ( .en(en), .clk(clk), .rst(rst), .q(c701ibus), .r(c701obus));
wire [temp_w*6-1:0] c702ibus;
wire [data_w*6-1:0] c702obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU702 ( .en(en), .clk(clk), .rst(rst), .q(c702ibus), .r(c702obus));
wire [temp_w*6-1:0] c703ibus;
wire [data_w*6-1:0] c703obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU703 ( .en(en), .clk(clk), .rst(rst), .q(c703ibus), .r(c703obus));
wire [temp_w*6-1:0] c704ibus;
wire [data_w*6-1:0] c704obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU704 ( .en(en), .clk(clk), .rst(rst), .q(c704ibus), .r(c704obus));
wire [temp_w*6-1:0] c705ibus;
wire [data_w*6-1:0] c705obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU705 ( .en(en), .clk(clk), .rst(rst), .q(c705ibus), .r(c705obus));
wire [temp_w*6-1:0] c706ibus;
wire [data_w*6-1:0] c706obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU706 ( .en(en), .clk(clk), .rst(rst), .q(c706ibus), .r(c706obus));
wire [temp_w*6-1:0] c707ibus;
wire [data_w*6-1:0] c707obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU707 ( .en(en), .clk(clk), .rst(rst), .q(c707ibus), .r(c707obus));
wire [temp_w*6-1:0] c708ibus;
wire [data_w*6-1:0] c708obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU708 ( .en(en), .clk(clk), .rst(rst), .q(c708ibus), .r(c708obus));
wire [temp_w*6-1:0] c709ibus;
wire [data_w*6-1:0] c709obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU709 ( .en(en), .clk(clk), .rst(rst), .q(c709ibus), .r(c709obus));
wire [temp_w*6-1:0] c710ibus;
wire [data_w*6-1:0] c710obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU710 ( .en(en), .clk(clk), .rst(rst), .q(c710ibus), .r(c710obus));
wire [temp_w*6-1:0] c711ibus;
wire [data_w*6-1:0] c711obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU711 ( .en(en), .clk(clk), .rst(rst), .q(c711ibus), .r(c711obus));
wire [temp_w*6-1:0] c712ibus;
wire [data_w*6-1:0] c712obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU712 ( .en(en), .clk(clk), .rst(rst), .q(c712ibus), .r(c712obus));
wire [temp_w*6-1:0] c713ibus;
wire [data_w*6-1:0] c713obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU713 ( .en(en), .clk(clk), .rst(rst), .q(c713ibus), .r(c713obus));
wire [temp_w*6-1:0] c714ibus;
wire [data_w*6-1:0] c714obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU714 ( .en(en), .clk(clk), .rst(rst), .q(c714ibus), .r(c714obus));
wire [temp_w*6-1:0] c715ibus;
wire [data_w*6-1:0] c715obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU715 ( .en(en), .clk(clk), .rst(rst), .q(c715ibus), .r(c715obus));
wire [temp_w*6-1:0] c716ibus;
wire [data_w*6-1:0] c716obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU716 ( .en(en), .clk(clk), .rst(rst), .q(c716ibus), .r(c716obus));
wire [temp_w*6-1:0] c717ibus;
wire [data_w*6-1:0] c717obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU717 ( .en(en), .clk(clk), .rst(rst), .q(c717ibus), .r(c717obus));
wire [temp_w*6-1:0] c718ibus;
wire [data_w*6-1:0] c718obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU718 ( .en(en), .clk(clk), .rst(rst), .q(c718ibus), .r(c718obus));
wire [temp_w*6-1:0] c719ibus;
wire [data_w*6-1:0] c719obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU719 ( .en(en), .clk(clk), .rst(rst), .q(c719ibus), .r(c719obus));
wire [temp_w*6-1:0] c720ibus;
wire [data_w*6-1:0] c720obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU720 ( .en(en), .clk(clk), .rst(rst), .q(c720ibus), .r(c720obus));
wire [temp_w*6-1:0] c721ibus;
wire [data_w*6-1:0] c721obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU721 ( .en(en), .clk(clk), .rst(rst), .q(c721ibus), .r(c721obus));
wire [temp_w*6-1:0] c722ibus;
wire [data_w*6-1:0] c722obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU722 ( .en(en), .clk(clk), .rst(rst), .q(c722ibus), .r(c722obus));
wire [temp_w*6-1:0] c723ibus;
wire [data_w*6-1:0] c723obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU723 ( .en(en), .clk(clk), .rst(rst), .q(c723ibus), .r(c723obus));
wire [temp_w*6-1:0] c724ibus;
wire [data_w*6-1:0] c724obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU724 ( .en(en), .clk(clk), .rst(rst), .q(c724ibus), .r(c724obus));
wire [temp_w*6-1:0] c725ibus;
wire [data_w*6-1:0] c725obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU725 ( .en(en), .clk(clk), .rst(rst), .q(c725ibus), .r(c725obus));
wire [temp_w*6-1:0] c726ibus;
wire [data_w*6-1:0] c726obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU726 ( .en(en), .clk(clk), .rst(rst), .q(c726ibus), .r(c726obus));
wire [temp_w*6-1:0] c727ibus;
wire [data_w*6-1:0] c727obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU727 ( .en(en), .clk(clk), .rst(rst), .q(c727ibus), .r(c727obus));
wire [temp_w*6-1:0] c728ibus;
wire [data_w*6-1:0] c728obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU728 ( .en(en), .clk(clk), .rst(rst), .q(c728ibus), .r(c728obus));
wire [temp_w*6-1:0] c729ibus;
wire [data_w*6-1:0] c729obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU729 ( .en(en), .clk(clk), .rst(rst), .q(c729ibus), .r(c729obus));
wire [temp_w*6-1:0] c730ibus;
wire [data_w*6-1:0] c730obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU730 ( .en(en), .clk(clk), .rst(rst), .q(c730ibus), .r(c730obus));
wire [temp_w*6-1:0] c731ibus;
wire [data_w*6-1:0] c731obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU731 ( .en(en), .clk(clk), .rst(rst), .q(c731ibus), .r(c731obus));
wire [temp_w*6-1:0] c732ibus;
wire [data_w*6-1:0] c732obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU732 ( .en(en), .clk(clk), .rst(rst), .q(c732ibus), .r(c732obus));
wire [temp_w*6-1:0] c733ibus;
wire [data_w*6-1:0] c733obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU733 ( .en(en), .clk(clk), .rst(rst), .q(c733ibus), .r(c733obus));
wire [temp_w*6-1:0] c734ibus;
wire [data_w*6-1:0] c734obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU734 ( .en(en), .clk(clk), .rst(rst), .q(c734ibus), .r(c734obus));
wire [temp_w*6-1:0] c735ibus;
wire [data_w*6-1:0] c735obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU735 ( .en(en), .clk(clk), .rst(rst), .q(c735ibus), .r(c735obus));
wire [temp_w*6-1:0] c736ibus;
wire [data_w*6-1:0] c736obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU736 ( .en(en), .clk(clk), .rst(rst), .q(c736ibus), .r(c736obus));
wire [temp_w*6-1:0] c737ibus;
wire [data_w*6-1:0] c737obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU737 ( .en(en), .clk(clk), .rst(rst), .q(c737ibus), .r(c737obus));
wire [temp_w*6-1:0] c738ibus;
wire [data_w*6-1:0] c738obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU738 ( .en(en), .clk(clk), .rst(rst), .q(c738ibus), .r(c738obus));
wire [temp_w*6-1:0] c739ibus;
wire [data_w*6-1:0] c739obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU739 ( .en(en), .clk(clk), .rst(rst), .q(c739ibus), .r(c739obus));
wire [temp_w*6-1:0] c740ibus;
wire [data_w*6-1:0] c740obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU740 ( .en(en), .clk(clk), .rst(rst), .q(c740ibus), .r(c740obus));
wire [temp_w*6-1:0] c741ibus;
wire [data_w*6-1:0] c741obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU741 ( .en(en), .clk(clk), .rst(rst), .q(c741ibus), .r(c741obus));
wire [temp_w*6-1:0] c742ibus;
wire [data_w*6-1:0] c742obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU742 ( .en(en), .clk(clk), .rst(rst), .q(c742ibus), .r(c742obus));
wire [temp_w*6-1:0] c743ibus;
wire [data_w*6-1:0] c743obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU743 ( .en(en), .clk(clk), .rst(rst), .q(c743ibus), .r(c743obus));
wire [temp_w*6-1:0] c744ibus;
wire [data_w*6-1:0] c744obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU744 ( .en(en), .clk(clk), .rst(rst), .q(c744ibus), .r(c744obus));
wire [temp_w*6-1:0] c745ibus;
wire [data_w*6-1:0] c745obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU745 ( .en(en), .clk(clk), .rst(rst), .q(c745ibus), .r(c745obus));
wire [temp_w*6-1:0] c746ibus;
wire [data_w*6-1:0] c746obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU746 ( .en(en), .clk(clk), .rst(rst), .q(c746ibus), .r(c746obus));
wire [temp_w*6-1:0] c747ibus;
wire [data_w*6-1:0] c747obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU747 ( .en(en), .clk(clk), .rst(rst), .q(c747ibus), .r(c747obus));
wire [temp_w*6-1:0] c748ibus;
wire [data_w*6-1:0] c748obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU748 ( .en(en), .clk(clk), .rst(rst), .q(c748ibus), .r(c748obus));
wire [temp_w*6-1:0] c749ibus;
wire [data_w*6-1:0] c749obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU749 ( .en(en), .clk(clk), .rst(rst), .q(c749ibus), .r(c749obus));
wire [temp_w*6-1:0] c750ibus;
wire [data_w*6-1:0] c750obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU750 ( .en(en), .clk(clk), .rst(rst), .q(c750ibus), .r(c750obus));
wire [temp_w*6-1:0] c751ibus;
wire [data_w*6-1:0] c751obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU751 ( .en(en), .clk(clk), .rst(rst), .q(c751ibus), .r(c751obus));
wire [temp_w*6-1:0] c752ibus;
wire [data_w*6-1:0] c752obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU752 ( .en(en), .clk(clk), .rst(rst), .q(c752ibus), .r(c752obus));
wire [temp_w*6-1:0] c753ibus;
wire [data_w*6-1:0] c753obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU753 ( .en(en), .clk(clk), .rst(rst), .q(c753ibus), .r(c753obus));
wire [temp_w*6-1:0] c754ibus;
wire [data_w*6-1:0] c754obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU754 ( .en(en), .clk(clk), .rst(rst), .q(c754ibus), .r(c754obus));
wire [temp_w*6-1:0] c755ibus;
wire [data_w*6-1:0] c755obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU755 ( .en(en), .clk(clk), .rst(rst), .q(c755ibus), .r(c755obus));
wire [temp_w*6-1:0] c756ibus;
wire [data_w*6-1:0] c756obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU756 ( .en(en), .clk(clk), .rst(rst), .q(c756ibus), .r(c756obus));
wire [temp_w*6-1:0] c757ibus;
wire [data_w*6-1:0] c757obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU757 ( .en(en), .clk(clk), .rst(rst), .q(c757ibus), .r(c757obus));
wire [temp_w*6-1:0] c758ibus;
wire [data_w*6-1:0] c758obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU758 ( .en(en), .clk(clk), .rst(rst), .q(c758ibus), .r(c758obus));
wire [temp_w*6-1:0] c759ibus;
wire [data_w*6-1:0] c759obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU759 ( .en(en), .clk(clk), .rst(rst), .q(c759ibus), .r(c759obus));
wire [temp_w*6-1:0] c760ibus;
wire [data_w*6-1:0] c760obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU760 ( .en(en), .clk(clk), .rst(rst), .q(c760ibus), .r(c760obus));
wire [temp_w*6-1:0] c761ibus;
wire [data_w*6-1:0] c761obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU761 ( .en(en), .clk(clk), .rst(rst), .q(c761ibus), .r(c761obus));
wire [temp_w*6-1:0] c762ibus;
wire [data_w*6-1:0] c762obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU762 ( .en(en), .clk(clk), .rst(rst), .q(c762ibus), .r(c762obus));
wire [temp_w*6-1:0] c763ibus;
wire [data_w*6-1:0] c763obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU763 ( .en(en), .clk(clk), .rst(rst), .q(c763ibus), .r(c763obus));
wire [temp_w*6-1:0] c764ibus;
wire [data_w*6-1:0] c764obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU764 ( .en(en), .clk(clk), .rst(rst), .q(c764ibus), .r(c764obus));
wire [temp_w*6-1:0] c765ibus;
wire [data_w*6-1:0] c765obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU765 ( .en(en), .clk(clk), .rst(rst), .q(c765ibus), .r(c765obus));
wire [temp_w*6-1:0] c766ibus;
wire [data_w*6-1:0] c766obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU766 ( .en(en), .clk(clk), .rst(rst), .q(c766ibus), .r(c766obus));
wire [temp_w*6-1:0] c767ibus;
wire [data_w*6-1:0] c767obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU767 ( .en(en), .clk(clk), .rst(rst), .q(c767ibus), .r(c767obus));
wire [temp_w*7-1:0] c768ibus;
wire [data_w*7-1:0] c768obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU768 ( .en(en), .clk(clk), .rst(rst), .q(c768ibus), .r(c768obus));
wire [temp_w*7-1:0] c769ibus;
wire [data_w*7-1:0] c769obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU769 ( .en(en), .clk(clk), .rst(rst), .q(c769ibus), .r(c769obus));
wire [temp_w*7-1:0] c770ibus;
wire [data_w*7-1:0] c770obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU770 ( .en(en), .clk(clk), .rst(rst), .q(c770ibus), .r(c770obus));
wire [temp_w*7-1:0] c771ibus;
wire [data_w*7-1:0] c771obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU771 ( .en(en), .clk(clk), .rst(rst), .q(c771ibus), .r(c771obus));
wire [temp_w*7-1:0] c772ibus;
wire [data_w*7-1:0] c772obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU772 ( .en(en), .clk(clk), .rst(rst), .q(c772ibus), .r(c772obus));
wire [temp_w*7-1:0] c773ibus;
wire [data_w*7-1:0] c773obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU773 ( .en(en), .clk(clk), .rst(rst), .q(c773ibus), .r(c773obus));
wire [temp_w*7-1:0] c774ibus;
wire [data_w*7-1:0] c774obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU774 ( .en(en), .clk(clk), .rst(rst), .q(c774ibus), .r(c774obus));
wire [temp_w*7-1:0] c775ibus;
wire [data_w*7-1:0] c775obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU775 ( .en(en), .clk(clk), .rst(rst), .q(c775ibus), .r(c775obus));
wire [temp_w*7-1:0] c776ibus;
wire [data_w*7-1:0] c776obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU776 ( .en(en), .clk(clk), .rst(rst), .q(c776ibus), .r(c776obus));
wire [temp_w*7-1:0] c777ibus;
wire [data_w*7-1:0] c777obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU777 ( .en(en), .clk(clk), .rst(rst), .q(c777ibus), .r(c777obus));
wire [temp_w*7-1:0] c778ibus;
wire [data_w*7-1:0] c778obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU778 ( .en(en), .clk(clk), .rst(rst), .q(c778ibus), .r(c778obus));
wire [temp_w*7-1:0] c779ibus;
wire [data_w*7-1:0] c779obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU779 ( .en(en), .clk(clk), .rst(rst), .q(c779ibus), .r(c779obus));
wire [temp_w*7-1:0] c780ibus;
wire [data_w*7-1:0] c780obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU780 ( .en(en), .clk(clk), .rst(rst), .q(c780ibus), .r(c780obus));
wire [temp_w*7-1:0] c781ibus;
wire [data_w*7-1:0] c781obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU781 ( .en(en), .clk(clk), .rst(rst), .q(c781ibus), .r(c781obus));
wire [temp_w*7-1:0] c782ibus;
wire [data_w*7-1:0] c782obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU782 ( .en(en), .clk(clk), .rst(rst), .q(c782ibus), .r(c782obus));
wire [temp_w*7-1:0] c783ibus;
wire [data_w*7-1:0] c783obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU783 ( .en(en), .clk(clk), .rst(rst), .q(c783ibus), .r(c783obus));
wire [temp_w*7-1:0] c784ibus;
wire [data_w*7-1:0] c784obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU784 ( .en(en), .clk(clk), .rst(rst), .q(c784ibus), .r(c784obus));
wire [temp_w*7-1:0] c785ibus;
wire [data_w*7-1:0] c785obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU785 ( .en(en), .clk(clk), .rst(rst), .q(c785ibus), .r(c785obus));
wire [temp_w*7-1:0] c786ibus;
wire [data_w*7-1:0] c786obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU786 ( .en(en), .clk(clk), .rst(rst), .q(c786ibus), .r(c786obus));
wire [temp_w*7-1:0] c787ibus;
wire [data_w*7-1:0] c787obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU787 ( .en(en), .clk(clk), .rst(rst), .q(c787ibus), .r(c787obus));
wire [temp_w*7-1:0] c788ibus;
wire [data_w*7-1:0] c788obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU788 ( .en(en), .clk(clk), .rst(rst), .q(c788ibus), .r(c788obus));
wire [temp_w*7-1:0] c789ibus;
wire [data_w*7-1:0] c789obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU789 ( .en(en), .clk(clk), .rst(rst), .q(c789ibus), .r(c789obus));
wire [temp_w*7-1:0] c790ibus;
wire [data_w*7-1:0] c790obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU790 ( .en(en), .clk(clk), .rst(rst), .q(c790ibus), .r(c790obus));
wire [temp_w*7-1:0] c791ibus;
wire [data_w*7-1:0] c791obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU791 ( .en(en), .clk(clk), .rst(rst), .q(c791ibus), .r(c791obus));
wire [temp_w*7-1:0] c792ibus;
wire [data_w*7-1:0] c792obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU792 ( .en(en), .clk(clk), .rst(rst), .q(c792ibus), .r(c792obus));
wire [temp_w*7-1:0] c793ibus;
wire [data_w*7-1:0] c793obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU793 ( .en(en), .clk(clk), .rst(rst), .q(c793ibus), .r(c793obus));
wire [temp_w*7-1:0] c794ibus;
wire [data_w*7-1:0] c794obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU794 ( .en(en), .clk(clk), .rst(rst), .q(c794ibus), .r(c794obus));
wire [temp_w*7-1:0] c795ibus;
wire [data_w*7-1:0] c795obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU795 ( .en(en), .clk(clk), .rst(rst), .q(c795ibus), .r(c795obus));
wire [temp_w*7-1:0] c796ibus;
wire [data_w*7-1:0] c796obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU796 ( .en(en), .clk(clk), .rst(rst), .q(c796ibus), .r(c796obus));
wire [temp_w*7-1:0] c797ibus;
wire [data_w*7-1:0] c797obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU797 ( .en(en), .clk(clk), .rst(rst), .q(c797ibus), .r(c797obus));
wire [temp_w*7-1:0] c798ibus;
wire [data_w*7-1:0] c798obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU798 ( .en(en), .clk(clk), .rst(rst), .q(c798ibus), .r(c798obus));
wire [temp_w*7-1:0] c799ibus;
wire [data_w*7-1:0] c799obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU799 ( .en(en), .clk(clk), .rst(rst), .q(c799ibus), .r(c799obus));
wire [temp_w*7-1:0] c800ibus;
wire [data_w*7-1:0] c800obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU800 ( .en(en), .clk(clk), .rst(rst), .q(c800ibus), .r(c800obus));
wire [temp_w*7-1:0] c801ibus;
wire [data_w*7-1:0] c801obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU801 ( .en(en), .clk(clk), .rst(rst), .q(c801ibus), .r(c801obus));
wire [temp_w*7-1:0] c802ibus;
wire [data_w*7-1:0] c802obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU802 ( .en(en), .clk(clk), .rst(rst), .q(c802ibus), .r(c802obus));
wire [temp_w*7-1:0] c803ibus;
wire [data_w*7-1:0] c803obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU803 ( .en(en), .clk(clk), .rst(rst), .q(c803ibus), .r(c803obus));
wire [temp_w*7-1:0] c804ibus;
wire [data_w*7-1:0] c804obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU804 ( .en(en), .clk(clk), .rst(rst), .q(c804ibus), .r(c804obus));
wire [temp_w*7-1:0] c805ibus;
wire [data_w*7-1:0] c805obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU805 ( .en(en), .clk(clk), .rst(rst), .q(c805ibus), .r(c805obus));
wire [temp_w*7-1:0] c806ibus;
wire [data_w*7-1:0] c806obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU806 ( .en(en), .clk(clk), .rst(rst), .q(c806ibus), .r(c806obus));
wire [temp_w*7-1:0] c807ibus;
wire [data_w*7-1:0] c807obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU807 ( .en(en), .clk(clk), .rst(rst), .q(c807ibus), .r(c807obus));
wire [temp_w*7-1:0] c808ibus;
wire [data_w*7-1:0] c808obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU808 ( .en(en), .clk(clk), .rst(rst), .q(c808ibus), .r(c808obus));
wire [temp_w*7-1:0] c809ibus;
wire [data_w*7-1:0] c809obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU809 ( .en(en), .clk(clk), .rst(rst), .q(c809ibus), .r(c809obus));
wire [temp_w*7-1:0] c810ibus;
wire [data_w*7-1:0] c810obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU810 ( .en(en), .clk(clk), .rst(rst), .q(c810ibus), .r(c810obus));
wire [temp_w*7-1:0] c811ibus;
wire [data_w*7-1:0] c811obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU811 ( .en(en), .clk(clk), .rst(rst), .q(c811ibus), .r(c811obus));
wire [temp_w*7-1:0] c812ibus;
wire [data_w*7-1:0] c812obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU812 ( .en(en), .clk(clk), .rst(rst), .q(c812ibus), .r(c812obus));
wire [temp_w*7-1:0] c813ibus;
wire [data_w*7-1:0] c813obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU813 ( .en(en), .clk(clk), .rst(rst), .q(c813ibus), .r(c813obus));
wire [temp_w*7-1:0] c814ibus;
wire [data_w*7-1:0] c814obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU814 ( .en(en), .clk(clk), .rst(rst), .q(c814ibus), .r(c814obus));
wire [temp_w*7-1:0] c815ibus;
wire [data_w*7-1:0] c815obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU815 ( .en(en), .clk(clk), .rst(rst), .q(c815ibus), .r(c815obus));
wire [temp_w*7-1:0] c816ibus;
wire [data_w*7-1:0] c816obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU816 ( .en(en), .clk(clk), .rst(rst), .q(c816ibus), .r(c816obus));
wire [temp_w*7-1:0] c817ibus;
wire [data_w*7-1:0] c817obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU817 ( .en(en), .clk(clk), .rst(rst), .q(c817ibus), .r(c817obus));
wire [temp_w*7-1:0] c818ibus;
wire [data_w*7-1:0] c818obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU818 ( .en(en), .clk(clk), .rst(rst), .q(c818ibus), .r(c818obus));
wire [temp_w*7-1:0] c819ibus;
wire [data_w*7-1:0] c819obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU819 ( .en(en), .clk(clk), .rst(rst), .q(c819ibus), .r(c819obus));
wire [temp_w*7-1:0] c820ibus;
wire [data_w*7-1:0] c820obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU820 ( .en(en), .clk(clk), .rst(rst), .q(c820ibus), .r(c820obus));
wire [temp_w*7-1:0] c821ibus;
wire [data_w*7-1:0] c821obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU821 ( .en(en), .clk(clk), .rst(rst), .q(c821ibus), .r(c821obus));
wire [temp_w*7-1:0] c822ibus;
wire [data_w*7-1:0] c822obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU822 ( .en(en), .clk(clk), .rst(rst), .q(c822ibus), .r(c822obus));
wire [temp_w*7-1:0] c823ibus;
wire [data_w*7-1:0] c823obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU823 ( .en(en), .clk(clk), .rst(rst), .q(c823ibus), .r(c823obus));
wire [temp_w*7-1:0] c824ibus;
wire [data_w*7-1:0] c824obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU824 ( .en(en), .clk(clk), .rst(rst), .q(c824ibus), .r(c824obus));
wire [temp_w*7-1:0] c825ibus;
wire [data_w*7-1:0] c825obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU825 ( .en(en), .clk(clk), .rst(rst), .q(c825ibus), .r(c825obus));
wire [temp_w*7-1:0] c826ibus;
wire [data_w*7-1:0] c826obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU826 ( .en(en), .clk(clk), .rst(rst), .q(c826ibus), .r(c826obus));
wire [temp_w*7-1:0] c827ibus;
wire [data_w*7-1:0] c827obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU827 ( .en(en), .clk(clk), .rst(rst), .q(c827ibus), .r(c827obus));
wire [temp_w*7-1:0] c828ibus;
wire [data_w*7-1:0] c828obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU828 ( .en(en), .clk(clk), .rst(rst), .q(c828ibus), .r(c828obus));
wire [temp_w*7-1:0] c829ibus;
wire [data_w*7-1:0] c829obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU829 ( .en(en), .clk(clk), .rst(rst), .q(c829ibus), .r(c829obus));
wire [temp_w*7-1:0] c830ibus;
wire [data_w*7-1:0] c830obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU830 ( .en(en), .clk(clk), .rst(rst), .q(c830ibus), .r(c830obus));
wire [temp_w*7-1:0] c831ibus;
wire [data_w*7-1:0] c831obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU831 ( .en(en), .clk(clk), .rst(rst), .q(c831ibus), .r(c831obus));
wire [temp_w*7-1:0] c832ibus;
wire [data_w*7-1:0] c832obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU832 ( .en(en), .clk(clk), .rst(rst), .q(c832ibus), .r(c832obus));
wire [temp_w*7-1:0] c833ibus;
wire [data_w*7-1:0] c833obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU833 ( .en(en), .clk(clk), .rst(rst), .q(c833ibus), .r(c833obus));
wire [temp_w*7-1:0] c834ibus;
wire [data_w*7-1:0] c834obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU834 ( .en(en), .clk(clk), .rst(rst), .q(c834ibus), .r(c834obus));
wire [temp_w*7-1:0] c835ibus;
wire [data_w*7-1:0] c835obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU835 ( .en(en), .clk(clk), .rst(rst), .q(c835ibus), .r(c835obus));
wire [temp_w*7-1:0] c836ibus;
wire [data_w*7-1:0] c836obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU836 ( .en(en), .clk(clk), .rst(rst), .q(c836ibus), .r(c836obus));
wire [temp_w*7-1:0] c837ibus;
wire [data_w*7-1:0] c837obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU837 ( .en(en), .clk(clk), .rst(rst), .q(c837ibus), .r(c837obus));
wire [temp_w*7-1:0] c838ibus;
wire [data_w*7-1:0] c838obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU838 ( .en(en), .clk(clk), .rst(rst), .q(c838ibus), .r(c838obus));
wire [temp_w*7-1:0] c839ibus;
wire [data_w*7-1:0] c839obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU839 ( .en(en), .clk(clk), .rst(rst), .q(c839ibus), .r(c839obus));
wire [temp_w*7-1:0] c840ibus;
wire [data_w*7-1:0] c840obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU840 ( .en(en), .clk(clk), .rst(rst), .q(c840ibus), .r(c840obus));
wire [temp_w*7-1:0] c841ibus;
wire [data_w*7-1:0] c841obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU841 ( .en(en), .clk(clk), .rst(rst), .q(c841ibus), .r(c841obus));
wire [temp_w*7-1:0] c842ibus;
wire [data_w*7-1:0] c842obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU842 ( .en(en), .clk(clk), .rst(rst), .q(c842ibus), .r(c842obus));
wire [temp_w*7-1:0] c843ibus;
wire [data_w*7-1:0] c843obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU843 ( .en(en), .clk(clk), .rst(rst), .q(c843ibus), .r(c843obus));
wire [temp_w*7-1:0] c844ibus;
wire [data_w*7-1:0] c844obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU844 ( .en(en), .clk(clk), .rst(rst), .q(c844ibus), .r(c844obus));
wire [temp_w*7-1:0] c845ibus;
wire [data_w*7-1:0] c845obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU845 ( .en(en), .clk(clk), .rst(rst), .q(c845ibus), .r(c845obus));
wire [temp_w*7-1:0] c846ibus;
wire [data_w*7-1:0] c846obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU846 ( .en(en), .clk(clk), .rst(rst), .q(c846ibus), .r(c846obus));
wire [temp_w*7-1:0] c847ibus;
wire [data_w*7-1:0] c847obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU847 ( .en(en), .clk(clk), .rst(rst), .q(c847ibus), .r(c847obus));
wire [temp_w*7-1:0] c848ibus;
wire [data_w*7-1:0] c848obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU848 ( .en(en), .clk(clk), .rst(rst), .q(c848ibus), .r(c848obus));
wire [temp_w*7-1:0] c849ibus;
wire [data_w*7-1:0] c849obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU849 ( .en(en), .clk(clk), .rst(rst), .q(c849ibus), .r(c849obus));
wire [temp_w*7-1:0] c850ibus;
wire [data_w*7-1:0] c850obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU850 ( .en(en), .clk(clk), .rst(rst), .q(c850ibus), .r(c850obus));
wire [temp_w*7-1:0] c851ibus;
wire [data_w*7-1:0] c851obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU851 ( .en(en), .clk(clk), .rst(rst), .q(c851ibus), .r(c851obus));
wire [temp_w*7-1:0] c852ibus;
wire [data_w*7-1:0] c852obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU852 ( .en(en), .clk(clk), .rst(rst), .q(c852ibus), .r(c852obus));
wire [temp_w*7-1:0] c853ibus;
wire [data_w*7-1:0] c853obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU853 ( .en(en), .clk(clk), .rst(rst), .q(c853ibus), .r(c853obus));
wire [temp_w*7-1:0] c854ibus;
wire [data_w*7-1:0] c854obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU854 ( .en(en), .clk(clk), .rst(rst), .q(c854ibus), .r(c854obus));
wire [temp_w*7-1:0] c855ibus;
wire [data_w*7-1:0] c855obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU855 ( .en(en), .clk(clk), .rst(rst), .q(c855ibus), .r(c855obus));
wire [temp_w*7-1:0] c856ibus;
wire [data_w*7-1:0] c856obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU856 ( .en(en), .clk(clk), .rst(rst), .q(c856ibus), .r(c856obus));
wire [temp_w*7-1:0] c857ibus;
wire [data_w*7-1:0] c857obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU857 ( .en(en), .clk(clk), .rst(rst), .q(c857ibus), .r(c857obus));
wire [temp_w*7-1:0] c858ibus;
wire [data_w*7-1:0] c858obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU858 ( .en(en), .clk(clk), .rst(rst), .q(c858ibus), .r(c858obus));
wire [temp_w*7-1:0] c859ibus;
wire [data_w*7-1:0] c859obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU859 ( .en(en), .clk(clk), .rst(rst), .q(c859ibus), .r(c859obus));
wire [temp_w*7-1:0] c860ibus;
wire [data_w*7-1:0] c860obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU860 ( .en(en), .clk(clk), .rst(rst), .q(c860ibus), .r(c860obus));
wire [temp_w*7-1:0] c861ibus;
wire [data_w*7-1:0] c861obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU861 ( .en(en), .clk(clk), .rst(rst), .q(c861ibus), .r(c861obus));
wire [temp_w*7-1:0] c862ibus;
wire [data_w*7-1:0] c862obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU862 ( .en(en), .clk(clk), .rst(rst), .q(c862ibus), .r(c862obus));
wire [temp_w*7-1:0] c863ibus;
wire [data_w*7-1:0] c863obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(7), .idx_w(idx_w)) CNU863 ( .en(en), .clk(clk), .rst(rst), .q(c863ibus), .r(c863obus));
wire [temp_w*6-1:0] c864ibus;
wire [data_w*6-1:0] c864obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU864 ( .en(en), .clk(clk), .rst(rst), .q(c864ibus), .r(c864obus));
wire [temp_w*6-1:0] c865ibus;
wire [data_w*6-1:0] c865obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU865 ( .en(en), .clk(clk), .rst(rst), .q(c865ibus), .r(c865obus));
wire [temp_w*6-1:0] c866ibus;
wire [data_w*6-1:0] c866obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU866 ( .en(en), .clk(clk), .rst(rst), .q(c866ibus), .r(c866obus));
wire [temp_w*6-1:0] c867ibus;
wire [data_w*6-1:0] c867obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU867 ( .en(en), .clk(clk), .rst(rst), .q(c867ibus), .r(c867obus));
wire [temp_w*6-1:0] c868ibus;
wire [data_w*6-1:0] c868obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU868 ( .en(en), .clk(clk), .rst(rst), .q(c868ibus), .r(c868obus));
wire [temp_w*6-1:0] c869ibus;
wire [data_w*6-1:0] c869obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU869 ( .en(en), .clk(clk), .rst(rst), .q(c869ibus), .r(c869obus));
wire [temp_w*6-1:0] c870ibus;
wire [data_w*6-1:0] c870obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU870 ( .en(en), .clk(clk), .rst(rst), .q(c870ibus), .r(c870obus));
wire [temp_w*6-1:0] c871ibus;
wire [data_w*6-1:0] c871obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU871 ( .en(en), .clk(clk), .rst(rst), .q(c871ibus), .r(c871obus));
wire [temp_w*6-1:0] c872ibus;
wire [data_w*6-1:0] c872obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU872 ( .en(en), .clk(clk), .rst(rst), .q(c872ibus), .r(c872obus));
wire [temp_w*6-1:0] c873ibus;
wire [data_w*6-1:0] c873obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU873 ( .en(en), .clk(clk), .rst(rst), .q(c873ibus), .r(c873obus));
wire [temp_w*6-1:0] c874ibus;
wire [data_w*6-1:0] c874obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU874 ( .en(en), .clk(clk), .rst(rst), .q(c874ibus), .r(c874obus));
wire [temp_w*6-1:0] c875ibus;
wire [data_w*6-1:0] c875obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU875 ( .en(en), .clk(clk), .rst(rst), .q(c875ibus), .r(c875obus));
wire [temp_w*6-1:0] c876ibus;
wire [data_w*6-1:0] c876obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU876 ( .en(en), .clk(clk), .rst(rst), .q(c876ibus), .r(c876obus));
wire [temp_w*6-1:0] c877ibus;
wire [data_w*6-1:0] c877obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU877 ( .en(en), .clk(clk), .rst(rst), .q(c877ibus), .r(c877obus));
wire [temp_w*6-1:0] c878ibus;
wire [data_w*6-1:0] c878obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU878 ( .en(en), .clk(clk), .rst(rst), .q(c878ibus), .r(c878obus));
wire [temp_w*6-1:0] c879ibus;
wire [data_w*6-1:0] c879obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU879 ( .en(en), .clk(clk), .rst(rst), .q(c879ibus), .r(c879obus));
wire [temp_w*6-1:0] c880ibus;
wire [data_w*6-1:0] c880obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU880 ( .en(en), .clk(clk), .rst(rst), .q(c880ibus), .r(c880obus));
wire [temp_w*6-1:0] c881ibus;
wire [data_w*6-1:0] c881obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU881 ( .en(en), .clk(clk), .rst(rst), .q(c881ibus), .r(c881obus));
wire [temp_w*6-1:0] c882ibus;
wire [data_w*6-1:0] c882obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU882 ( .en(en), .clk(clk), .rst(rst), .q(c882ibus), .r(c882obus));
wire [temp_w*6-1:0] c883ibus;
wire [data_w*6-1:0] c883obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU883 ( .en(en), .clk(clk), .rst(rst), .q(c883ibus), .r(c883obus));
wire [temp_w*6-1:0] c884ibus;
wire [data_w*6-1:0] c884obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU884 ( .en(en), .clk(clk), .rst(rst), .q(c884ibus), .r(c884obus));
wire [temp_w*6-1:0] c885ibus;
wire [data_w*6-1:0] c885obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU885 ( .en(en), .clk(clk), .rst(rst), .q(c885ibus), .r(c885obus));
wire [temp_w*6-1:0] c886ibus;
wire [data_w*6-1:0] c886obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU886 ( .en(en), .clk(clk), .rst(rst), .q(c886ibus), .r(c886obus));
wire [temp_w*6-1:0] c887ibus;
wire [data_w*6-1:0] c887obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU887 ( .en(en), .clk(clk), .rst(rst), .q(c887ibus), .r(c887obus));
wire [temp_w*6-1:0] c888ibus;
wire [data_w*6-1:0] c888obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU888 ( .en(en), .clk(clk), .rst(rst), .q(c888ibus), .r(c888obus));
wire [temp_w*6-1:0] c889ibus;
wire [data_w*6-1:0] c889obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU889 ( .en(en), .clk(clk), .rst(rst), .q(c889ibus), .r(c889obus));
wire [temp_w*6-1:0] c890ibus;
wire [data_w*6-1:0] c890obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU890 ( .en(en), .clk(clk), .rst(rst), .q(c890ibus), .r(c890obus));
wire [temp_w*6-1:0] c891ibus;
wire [data_w*6-1:0] c891obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU891 ( .en(en), .clk(clk), .rst(rst), .q(c891ibus), .r(c891obus));
wire [temp_w*6-1:0] c892ibus;
wire [data_w*6-1:0] c892obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU892 ( .en(en), .clk(clk), .rst(rst), .q(c892ibus), .r(c892obus));
wire [temp_w*6-1:0] c893ibus;
wire [data_w*6-1:0] c893obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU893 ( .en(en), .clk(clk), .rst(rst), .q(c893ibus), .r(c893obus));
wire [temp_w*6-1:0] c894ibus;
wire [data_w*6-1:0] c894obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU894 ( .en(en), .clk(clk), .rst(rst), .q(c894ibus), .r(c894obus));
wire [temp_w*6-1:0] c895ibus;
wire [data_w*6-1:0] c895obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU895 ( .en(en), .clk(clk), .rst(rst), .q(c895ibus), .r(c895obus));
wire [temp_w*6-1:0] c896ibus;
wire [data_w*6-1:0] c896obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU896 ( .en(en), .clk(clk), .rst(rst), .q(c896ibus), .r(c896obus));
wire [temp_w*6-1:0] c897ibus;
wire [data_w*6-1:0] c897obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU897 ( .en(en), .clk(clk), .rst(rst), .q(c897ibus), .r(c897obus));
wire [temp_w*6-1:0] c898ibus;
wire [data_w*6-1:0] c898obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU898 ( .en(en), .clk(clk), .rst(rst), .q(c898ibus), .r(c898obus));
wire [temp_w*6-1:0] c899ibus;
wire [data_w*6-1:0] c899obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU899 ( .en(en), .clk(clk), .rst(rst), .q(c899ibus), .r(c899obus));
wire [temp_w*6-1:0] c900ibus;
wire [data_w*6-1:0] c900obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU900 ( .en(en), .clk(clk), .rst(rst), .q(c900ibus), .r(c900obus));
wire [temp_w*6-1:0] c901ibus;
wire [data_w*6-1:0] c901obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU901 ( .en(en), .clk(clk), .rst(rst), .q(c901ibus), .r(c901obus));
wire [temp_w*6-1:0] c902ibus;
wire [data_w*6-1:0] c902obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU902 ( .en(en), .clk(clk), .rst(rst), .q(c902ibus), .r(c902obus));
wire [temp_w*6-1:0] c903ibus;
wire [data_w*6-1:0] c903obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU903 ( .en(en), .clk(clk), .rst(rst), .q(c903ibus), .r(c903obus));
wire [temp_w*6-1:0] c904ibus;
wire [data_w*6-1:0] c904obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU904 ( .en(en), .clk(clk), .rst(rst), .q(c904ibus), .r(c904obus));
wire [temp_w*6-1:0] c905ibus;
wire [data_w*6-1:0] c905obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU905 ( .en(en), .clk(clk), .rst(rst), .q(c905ibus), .r(c905obus));
wire [temp_w*6-1:0] c906ibus;
wire [data_w*6-1:0] c906obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU906 ( .en(en), .clk(clk), .rst(rst), .q(c906ibus), .r(c906obus));
wire [temp_w*6-1:0] c907ibus;
wire [data_w*6-1:0] c907obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU907 ( .en(en), .clk(clk), .rst(rst), .q(c907ibus), .r(c907obus));
wire [temp_w*6-1:0] c908ibus;
wire [data_w*6-1:0] c908obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU908 ( .en(en), .clk(clk), .rst(rst), .q(c908ibus), .r(c908obus));
wire [temp_w*6-1:0] c909ibus;
wire [data_w*6-1:0] c909obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU909 ( .en(en), .clk(clk), .rst(rst), .q(c909ibus), .r(c909obus));
wire [temp_w*6-1:0] c910ibus;
wire [data_w*6-1:0] c910obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU910 ( .en(en), .clk(clk), .rst(rst), .q(c910ibus), .r(c910obus));
wire [temp_w*6-1:0] c911ibus;
wire [data_w*6-1:0] c911obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU911 ( .en(en), .clk(clk), .rst(rst), .q(c911ibus), .r(c911obus));
wire [temp_w*6-1:0] c912ibus;
wire [data_w*6-1:0] c912obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU912 ( .en(en), .clk(clk), .rst(rst), .q(c912ibus), .r(c912obus));
wire [temp_w*6-1:0] c913ibus;
wire [data_w*6-1:0] c913obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU913 ( .en(en), .clk(clk), .rst(rst), .q(c913ibus), .r(c913obus));
wire [temp_w*6-1:0] c914ibus;
wire [data_w*6-1:0] c914obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU914 ( .en(en), .clk(clk), .rst(rst), .q(c914ibus), .r(c914obus));
wire [temp_w*6-1:0] c915ibus;
wire [data_w*6-1:0] c915obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU915 ( .en(en), .clk(clk), .rst(rst), .q(c915ibus), .r(c915obus));
wire [temp_w*6-1:0] c916ibus;
wire [data_w*6-1:0] c916obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU916 ( .en(en), .clk(clk), .rst(rst), .q(c916ibus), .r(c916obus));
wire [temp_w*6-1:0] c917ibus;
wire [data_w*6-1:0] c917obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU917 ( .en(en), .clk(clk), .rst(rst), .q(c917ibus), .r(c917obus));
wire [temp_w*6-1:0] c918ibus;
wire [data_w*6-1:0] c918obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU918 ( .en(en), .clk(clk), .rst(rst), .q(c918ibus), .r(c918obus));
wire [temp_w*6-1:0] c919ibus;
wire [data_w*6-1:0] c919obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU919 ( .en(en), .clk(clk), .rst(rst), .q(c919ibus), .r(c919obus));
wire [temp_w*6-1:0] c920ibus;
wire [data_w*6-1:0] c920obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU920 ( .en(en), .clk(clk), .rst(rst), .q(c920ibus), .r(c920obus));
wire [temp_w*6-1:0] c921ibus;
wire [data_w*6-1:0] c921obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU921 ( .en(en), .clk(clk), .rst(rst), .q(c921ibus), .r(c921obus));
wire [temp_w*6-1:0] c922ibus;
wire [data_w*6-1:0] c922obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU922 ( .en(en), .clk(clk), .rst(rst), .q(c922ibus), .r(c922obus));
wire [temp_w*6-1:0] c923ibus;
wire [data_w*6-1:0] c923obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU923 ( .en(en), .clk(clk), .rst(rst), .q(c923ibus), .r(c923obus));
wire [temp_w*6-1:0] c924ibus;
wire [data_w*6-1:0] c924obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU924 ( .en(en), .clk(clk), .rst(rst), .q(c924ibus), .r(c924obus));
wire [temp_w*6-1:0] c925ibus;
wire [data_w*6-1:0] c925obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU925 ( .en(en), .clk(clk), .rst(rst), .q(c925ibus), .r(c925obus));
wire [temp_w*6-1:0] c926ibus;
wire [data_w*6-1:0] c926obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU926 ( .en(en), .clk(clk), .rst(rst), .q(c926ibus), .r(c926obus));
wire [temp_w*6-1:0] c927ibus;
wire [data_w*6-1:0] c927obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU927 ( .en(en), .clk(clk), .rst(rst), .q(c927ibus), .r(c927obus));
wire [temp_w*6-1:0] c928ibus;
wire [data_w*6-1:0] c928obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU928 ( .en(en), .clk(clk), .rst(rst), .q(c928ibus), .r(c928obus));
wire [temp_w*6-1:0] c929ibus;
wire [data_w*6-1:0] c929obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU929 ( .en(en), .clk(clk), .rst(rst), .q(c929ibus), .r(c929obus));
wire [temp_w*6-1:0] c930ibus;
wire [data_w*6-1:0] c930obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU930 ( .en(en), .clk(clk), .rst(rst), .q(c930ibus), .r(c930obus));
wire [temp_w*6-1:0] c931ibus;
wire [data_w*6-1:0] c931obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU931 ( .en(en), .clk(clk), .rst(rst), .q(c931ibus), .r(c931obus));
wire [temp_w*6-1:0] c932ibus;
wire [data_w*6-1:0] c932obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU932 ( .en(en), .clk(clk), .rst(rst), .q(c932ibus), .r(c932obus));
wire [temp_w*6-1:0] c933ibus;
wire [data_w*6-1:0] c933obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU933 ( .en(en), .clk(clk), .rst(rst), .q(c933ibus), .r(c933obus));
wire [temp_w*6-1:0] c934ibus;
wire [data_w*6-1:0] c934obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU934 ( .en(en), .clk(clk), .rst(rst), .q(c934ibus), .r(c934obus));
wire [temp_w*6-1:0] c935ibus;
wire [data_w*6-1:0] c935obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU935 ( .en(en), .clk(clk), .rst(rst), .q(c935ibus), .r(c935obus));
wire [temp_w*6-1:0] c936ibus;
wire [data_w*6-1:0] c936obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU936 ( .en(en), .clk(clk), .rst(rst), .q(c936ibus), .r(c936obus));
wire [temp_w*6-1:0] c937ibus;
wire [data_w*6-1:0] c937obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU937 ( .en(en), .clk(clk), .rst(rst), .q(c937ibus), .r(c937obus));
wire [temp_w*6-1:0] c938ibus;
wire [data_w*6-1:0] c938obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU938 ( .en(en), .clk(clk), .rst(rst), .q(c938ibus), .r(c938obus));
wire [temp_w*6-1:0] c939ibus;
wire [data_w*6-1:0] c939obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU939 ( .en(en), .clk(clk), .rst(rst), .q(c939ibus), .r(c939obus));
wire [temp_w*6-1:0] c940ibus;
wire [data_w*6-1:0] c940obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU940 ( .en(en), .clk(clk), .rst(rst), .q(c940ibus), .r(c940obus));
wire [temp_w*6-1:0] c941ibus;
wire [data_w*6-1:0] c941obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU941 ( .en(en), .clk(clk), .rst(rst), .q(c941ibus), .r(c941obus));
wire [temp_w*6-1:0] c942ibus;
wire [data_w*6-1:0] c942obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU942 ( .en(en), .clk(clk), .rst(rst), .q(c942ibus), .r(c942obus));
wire [temp_w*6-1:0] c943ibus;
wire [data_w*6-1:0] c943obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU943 ( .en(en), .clk(clk), .rst(rst), .q(c943ibus), .r(c943obus));
wire [temp_w*6-1:0] c944ibus;
wire [data_w*6-1:0] c944obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU944 ( .en(en), .clk(clk), .rst(rst), .q(c944ibus), .r(c944obus));
wire [temp_w*6-1:0] c945ibus;
wire [data_w*6-1:0] c945obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU945 ( .en(en), .clk(clk), .rst(rst), .q(c945ibus), .r(c945obus));
wire [temp_w*6-1:0] c946ibus;
wire [data_w*6-1:0] c946obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU946 ( .en(en), .clk(clk), .rst(rst), .q(c946ibus), .r(c946obus));
wire [temp_w*6-1:0] c947ibus;
wire [data_w*6-1:0] c947obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU947 ( .en(en), .clk(clk), .rst(rst), .q(c947ibus), .r(c947obus));
wire [temp_w*6-1:0] c948ibus;
wire [data_w*6-1:0] c948obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU948 ( .en(en), .clk(clk), .rst(rst), .q(c948ibus), .r(c948obus));
wire [temp_w*6-1:0] c949ibus;
wire [data_w*6-1:0] c949obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU949 ( .en(en), .clk(clk), .rst(rst), .q(c949ibus), .r(c949obus));
wire [temp_w*6-1:0] c950ibus;
wire [data_w*6-1:0] c950obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU950 ( .en(en), .clk(clk), .rst(rst), .q(c950ibus), .r(c950obus));
wire [temp_w*6-1:0] c951ibus;
wire [data_w*6-1:0] c951obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU951 ( .en(en), .clk(clk), .rst(rst), .q(c951ibus), .r(c951obus));
wire [temp_w*6-1:0] c952ibus;
wire [data_w*6-1:0] c952obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU952 ( .en(en), .clk(clk), .rst(rst), .q(c952ibus), .r(c952obus));
wire [temp_w*6-1:0] c953ibus;
wire [data_w*6-1:0] c953obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU953 ( .en(en), .clk(clk), .rst(rst), .q(c953ibus), .r(c953obus));
wire [temp_w*6-1:0] c954ibus;
wire [data_w*6-1:0] c954obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU954 ( .en(en), .clk(clk), .rst(rst), .q(c954ibus), .r(c954obus));
wire [temp_w*6-1:0] c955ibus;
wire [data_w*6-1:0] c955obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU955 ( .en(en), .clk(clk), .rst(rst), .q(c955ibus), .r(c955obus));
wire [temp_w*6-1:0] c956ibus;
wire [data_w*6-1:0] c956obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU956 ( .en(en), .clk(clk), .rst(rst), .q(c956ibus), .r(c956obus));
wire [temp_w*6-1:0] c957ibus;
wire [data_w*6-1:0] c957obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU957 ( .en(en), .clk(clk), .rst(rst), .q(c957ibus), .r(c957obus));
wire [temp_w*6-1:0] c958ibus;
wire [data_w*6-1:0] c958obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU958 ( .en(en), .clk(clk), .rst(rst), .q(c958ibus), .r(c958obus));
wire [temp_w*6-1:0] c959ibus;
wire [data_w*6-1:0] c959obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU959 ( .en(en), .clk(clk), .rst(rst), .q(c959ibus), .r(c959obus));
wire [temp_w*6-1:0] c960ibus;
wire [data_w*6-1:0] c960obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU960 ( .en(en), .clk(clk), .rst(rst), .q(c960ibus), .r(c960obus));
wire [temp_w*6-1:0] c961ibus;
wire [data_w*6-1:0] c961obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU961 ( .en(en), .clk(clk), .rst(rst), .q(c961ibus), .r(c961obus));
wire [temp_w*6-1:0] c962ibus;
wire [data_w*6-1:0] c962obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU962 ( .en(en), .clk(clk), .rst(rst), .q(c962ibus), .r(c962obus));
wire [temp_w*6-1:0] c963ibus;
wire [data_w*6-1:0] c963obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU963 ( .en(en), .clk(clk), .rst(rst), .q(c963ibus), .r(c963obus));
wire [temp_w*6-1:0] c964ibus;
wire [data_w*6-1:0] c964obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU964 ( .en(en), .clk(clk), .rst(rst), .q(c964ibus), .r(c964obus));
wire [temp_w*6-1:0] c965ibus;
wire [data_w*6-1:0] c965obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU965 ( .en(en), .clk(clk), .rst(rst), .q(c965ibus), .r(c965obus));
wire [temp_w*6-1:0] c966ibus;
wire [data_w*6-1:0] c966obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU966 ( .en(en), .clk(clk), .rst(rst), .q(c966ibus), .r(c966obus));
wire [temp_w*6-1:0] c967ibus;
wire [data_w*6-1:0] c967obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU967 ( .en(en), .clk(clk), .rst(rst), .q(c967ibus), .r(c967obus));
wire [temp_w*6-1:0] c968ibus;
wire [data_w*6-1:0] c968obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU968 ( .en(en), .clk(clk), .rst(rst), .q(c968ibus), .r(c968obus));
wire [temp_w*6-1:0] c969ibus;
wire [data_w*6-1:0] c969obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU969 ( .en(en), .clk(clk), .rst(rst), .q(c969ibus), .r(c969obus));
wire [temp_w*6-1:0] c970ibus;
wire [data_w*6-1:0] c970obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU970 ( .en(en), .clk(clk), .rst(rst), .q(c970ibus), .r(c970obus));
wire [temp_w*6-1:0] c971ibus;
wire [data_w*6-1:0] c971obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU971 ( .en(en), .clk(clk), .rst(rst), .q(c971ibus), .r(c971obus));
wire [temp_w*6-1:0] c972ibus;
wire [data_w*6-1:0] c972obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU972 ( .en(en), .clk(clk), .rst(rst), .q(c972ibus), .r(c972obus));
wire [temp_w*6-1:0] c973ibus;
wire [data_w*6-1:0] c973obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU973 ( .en(en), .clk(clk), .rst(rst), .q(c973ibus), .r(c973obus));
wire [temp_w*6-1:0] c974ibus;
wire [data_w*6-1:0] c974obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU974 ( .en(en), .clk(clk), .rst(rst), .q(c974ibus), .r(c974obus));
wire [temp_w*6-1:0] c975ibus;
wire [data_w*6-1:0] c975obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU975 ( .en(en), .clk(clk), .rst(rst), .q(c975ibus), .r(c975obus));
wire [temp_w*6-1:0] c976ibus;
wire [data_w*6-1:0] c976obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU976 ( .en(en), .clk(clk), .rst(rst), .q(c976ibus), .r(c976obus));
wire [temp_w*6-1:0] c977ibus;
wire [data_w*6-1:0] c977obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU977 ( .en(en), .clk(clk), .rst(rst), .q(c977ibus), .r(c977obus));
wire [temp_w*6-1:0] c978ibus;
wire [data_w*6-1:0] c978obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU978 ( .en(en), .clk(clk), .rst(rst), .q(c978ibus), .r(c978obus));
wire [temp_w*6-1:0] c979ibus;
wire [data_w*6-1:0] c979obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU979 ( .en(en), .clk(clk), .rst(rst), .q(c979ibus), .r(c979obus));
wire [temp_w*6-1:0] c980ibus;
wire [data_w*6-1:0] c980obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU980 ( .en(en), .clk(clk), .rst(rst), .q(c980ibus), .r(c980obus));
wire [temp_w*6-1:0] c981ibus;
wire [data_w*6-1:0] c981obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU981 ( .en(en), .clk(clk), .rst(rst), .q(c981ibus), .r(c981obus));
wire [temp_w*6-1:0] c982ibus;
wire [data_w*6-1:0] c982obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU982 ( .en(en), .clk(clk), .rst(rst), .q(c982ibus), .r(c982obus));
wire [temp_w*6-1:0] c983ibus;
wire [data_w*6-1:0] c983obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU983 ( .en(en), .clk(clk), .rst(rst), .q(c983ibus), .r(c983obus));
wire [temp_w*6-1:0] c984ibus;
wire [data_w*6-1:0] c984obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU984 ( .en(en), .clk(clk), .rst(rst), .q(c984ibus), .r(c984obus));
wire [temp_w*6-1:0] c985ibus;
wire [data_w*6-1:0] c985obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU985 ( .en(en), .clk(clk), .rst(rst), .q(c985ibus), .r(c985obus));
wire [temp_w*6-1:0] c986ibus;
wire [data_w*6-1:0] c986obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU986 ( .en(en), .clk(clk), .rst(rst), .q(c986ibus), .r(c986obus));
wire [temp_w*6-1:0] c987ibus;
wire [data_w*6-1:0] c987obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU987 ( .en(en), .clk(clk), .rst(rst), .q(c987ibus), .r(c987obus));
wire [temp_w*6-1:0] c988ibus;
wire [data_w*6-1:0] c988obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU988 ( .en(en), .clk(clk), .rst(rst), .q(c988ibus), .r(c988obus));
wire [temp_w*6-1:0] c989ibus;
wire [data_w*6-1:0] c989obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU989 ( .en(en), .clk(clk), .rst(rst), .q(c989ibus), .r(c989obus));
wire [temp_w*6-1:0] c990ibus;
wire [data_w*6-1:0] c990obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU990 ( .en(en), .clk(clk), .rst(rst), .q(c990ibus), .r(c990obus));
wire [temp_w*6-1:0] c991ibus;
wire [data_w*6-1:0] c991obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU991 ( .en(en), .clk(clk), .rst(rst), .q(c991ibus), .r(c991obus));
wire [temp_w*6-1:0] c992ibus;
wire [data_w*6-1:0] c992obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU992 ( .en(en), .clk(clk), .rst(rst), .q(c992ibus), .r(c992obus));
wire [temp_w*6-1:0] c993ibus;
wire [data_w*6-1:0] c993obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU993 ( .en(en), .clk(clk), .rst(rst), .q(c993ibus), .r(c993obus));
wire [temp_w*6-1:0] c994ibus;
wire [data_w*6-1:0] c994obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU994 ( .en(en), .clk(clk), .rst(rst), .q(c994ibus), .r(c994obus));
wire [temp_w*6-1:0] c995ibus;
wire [data_w*6-1:0] c995obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU995 ( .en(en), .clk(clk), .rst(rst), .q(c995ibus), .r(c995obus));
wire [temp_w*6-1:0] c996ibus;
wire [data_w*6-1:0] c996obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU996 ( .en(en), .clk(clk), .rst(rst), .q(c996ibus), .r(c996obus));
wire [temp_w*6-1:0] c997ibus;
wire [data_w*6-1:0] c997obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU997 ( .en(en), .clk(clk), .rst(rst), .q(c997ibus), .r(c997obus));
wire [temp_w*6-1:0] c998ibus;
wire [data_w*6-1:0] c998obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU998 ( .en(en), .clk(clk), .rst(rst), .q(c998ibus), .r(c998obus));
wire [temp_w*6-1:0] c999ibus;
wire [data_w*6-1:0] c999obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU999 ( .en(en), .clk(clk), .rst(rst), .q(c999ibus), .r(c999obus));
wire [temp_w*6-1:0] c1000ibus;
wire [data_w*6-1:0] c1000obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1000 ( .en(en), .clk(clk), .rst(rst), .q(c1000ibus), .r(c1000obus));
wire [temp_w*6-1:0] c1001ibus;
wire [data_w*6-1:0] c1001obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1001 ( .en(en), .clk(clk), .rst(rst), .q(c1001ibus), .r(c1001obus));
wire [temp_w*6-1:0] c1002ibus;
wire [data_w*6-1:0] c1002obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1002 ( .en(en), .clk(clk), .rst(rst), .q(c1002ibus), .r(c1002obus));
wire [temp_w*6-1:0] c1003ibus;
wire [data_w*6-1:0] c1003obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1003 ( .en(en), .clk(clk), .rst(rst), .q(c1003ibus), .r(c1003obus));
wire [temp_w*6-1:0] c1004ibus;
wire [data_w*6-1:0] c1004obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1004 ( .en(en), .clk(clk), .rst(rst), .q(c1004ibus), .r(c1004obus));
wire [temp_w*6-1:0] c1005ibus;
wire [data_w*6-1:0] c1005obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1005 ( .en(en), .clk(clk), .rst(rst), .q(c1005ibus), .r(c1005obus));
wire [temp_w*6-1:0] c1006ibus;
wire [data_w*6-1:0] c1006obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1006 ( .en(en), .clk(clk), .rst(rst), .q(c1006ibus), .r(c1006obus));
wire [temp_w*6-1:0] c1007ibus;
wire [data_w*6-1:0] c1007obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1007 ( .en(en), .clk(clk), .rst(rst), .q(c1007ibus), .r(c1007obus));
wire [temp_w*6-1:0] c1008ibus;
wire [data_w*6-1:0] c1008obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1008 ( .en(en), .clk(clk), .rst(rst), .q(c1008ibus), .r(c1008obus));
wire [temp_w*6-1:0] c1009ibus;
wire [data_w*6-1:0] c1009obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1009 ( .en(en), .clk(clk), .rst(rst), .q(c1009ibus), .r(c1009obus));
wire [temp_w*6-1:0] c1010ibus;
wire [data_w*6-1:0] c1010obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1010 ( .en(en), .clk(clk), .rst(rst), .q(c1010ibus), .r(c1010obus));
wire [temp_w*6-1:0] c1011ibus;
wire [data_w*6-1:0] c1011obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1011 ( .en(en), .clk(clk), .rst(rst), .q(c1011ibus), .r(c1011obus));
wire [temp_w*6-1:0] c1012ibus;
wire [data_w*6-1:0] c1012obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1012 ( .en(en), .clk(clk), .rst(rst), .q(c1012ibus), .r(c1012obus));
wire [temp_w*6-1:0] c1013ibus;
wire [data_w*6-1:0] c1013obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1013 ( .en(en), .clk(clk), .rst(rst), .q(c1013ibus), .r(c1013obus));
wire [temp_w*6-1:0] c1014ibus;
wire [data_w*6-1:0] c1014obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1014 ( .en(en), .clk(clk), .rst(rst), .q(c1014ibus), .r(c1014obus));
wire [temp_w*6-1:0] c1015ibus;
wire [data_w*6-1:0] c1015obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1015 ( .en(en), .clk(clk), .rst(rst), .q(c1015ibus), .r(c1015obus));
wire [temp_w*6-1:0] c1016ibus;
wire [data_w*6-1:0] c1016obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1016 ( .en(en), .clk(clk), .rst(rst), .q(c1016ibus), .r(c1016obus));
wire [temp_w*6-1:0] c1017ibus;
wire [data_w*6-1:0] c1017obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1017 ( .en(en), .clk(clk), .rst(rst), .q(c1017ibus), .r(c1017obus));
wire [temp_w*6-1:0] c1018ibus;
wire [data_w*6-1:0] c1018obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1018 ( .en(en), .clk(clk), .rst(rst), .q(c1018ibus), .r(c1018obus));
wire [temp_w*6-1:0] c1019ibus;
wire [data_w*6-1:0] c1019obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1019 ( .en(en), .clk(clk), .rst(rst), .q(c1019ibus), .r(c1019obus));
wire [temp_w*6-1:0] c1020ibus;
wire [data_w*6-1:0] c1020obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1020 ( .en(en), .clk(clk), .rst(rst), .q(c1020ibus), .r(c1020obus));
wire [temp_w*6-1:0] c1021ibus;
wire [data_w*6-1:0] c1021obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1021 ( .en(en), .clk(clk), .rst(rst), .q(c1021ibus), .r(c1021obus));
wire [temp_w*6-1:0] c1022ibus;
wire [data_w*6-1:0] c1022obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1022 ( .en(en), .clk(clk), .rst(rst), .q(c1022ibus), .r(c1022obus));
wire [temp_w*6-1:0] c1023ibus;
wire [data_w*6-1:0] c1023obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1023 ( .en(en), .clk(clk), .rst(rst), .q(c1023ibus), .r(c1023obus));
wire [temp_w*6-1:0] c1024ibus;
wire [data_w*6-1:0] c1024obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1024 ( .en(en), .clk(clk), .rst(rst), .q(c1024ibus), .r(c1024obus));
wire [temp_w*6-1:0] c1025ibus;
wire [data_w*6-1:0] c1025obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1025 ( .en(en), .clk(clk), .rst(rst), .q(c1025ibus), .r(c1025obus));
wire [temp_w*6-1:0] c1026ibus;
wire [data_w*6-1:0] c1026obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1026 ( .en(en), .clk(clk), .rst(rst), .q(c1026ibus), .r(c1026obus));
wire [temp_w*6-1:0] c1027ibus;
wire [data_w*6-1:0] c1027obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1027 ( .en(en), .clk(clk), .rst(rst), .q(c1027ibus), .r(c1027obus));
wire [temp_w*6-1:0] c1028ibus;
wire [data_w*6-1:0] c1028obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1028 ( .en(en), .clk(clk), .rst(rst), .q(c1028ibus), .r(c1028obus));
wire [temp_w*6-1:0] c1029ibus;
wire [data_w*6-1:0] c1029obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1029 ( .en(en), .clk(clk), .rst(rst), .q(c1029ibus), .r(c1029obus));
wire [temp_w*6-1:0] c1030ibus;
wire [data_w*6-1:0] c1030obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1030 ( .en(en), .clk(clk), .rst(rst), .q(c1030ibus), .r(c1030obus));
wire [temp_w*6-1:0] c1031ibus;
wire [data_w*6-1:0] c1031obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1031 ( .en(en), .clk(clk), .rst(rst), .q(c1031ibus), .r(c1031obus));
wire [temp_w*6-1:0] c1032ibus;
wire [data_w*6-1:0] c1032obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1032 ( .en(en), .clk(clk), .rst(rst), .q(c1032ibus), .r(c1032obus));
wire [temp_w*6-1:0] c1033ibus;
wire [data_w*6-1:0] c1033obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1033 ( .en(en), .clk(clk), .rst(rst), .q(c1033ibus), .r(c1033obus));
wire [temp_w*6-1:0] c1034ibus;
wire [data_w*6-1:0] c1034obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1034 ( .en(en), .clk(clk), .rst(rst), .q(c1034ibus), .r(c1034obus));
wire [temp_w*6-1:0] c1035ibus;
wire [data_w*6-1:0] c1035obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1035 ( .en(en), .clk(clk), .rst(rst), .q(c1035ibus), .r(c1035obus));
wire [temp_w*6-1:0] c1036ibus;
wire [data_w*6-1:0] c1036obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1036 ( .en(en), .clk(clk), .rst(rst), .q(c1036ibus), .r(c1036obus));
wire [temp_w*6-1:0] c1037ibus;
wire [data_w*6-1:0] c1037obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1037 ( .en(en), .clk(clk), .rst(rst), .q(c1037ibus), .r(c1037obus));
wire [temp_w*6-1:0] c1038ibus;
wire [data_w*6-1:0] c1038obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1038 ( .en(en), .clk(clk), .rst(rst), .q(c1038ibus), .r(c1038obus));
wire [temp_w*6-1:0] c1039ibus;
wire [data_w*6-1:0] c1039obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1039 ( .en(en), .clk(clk), .rst(rst), .q(c1039ibus), .r(c1039obus));
wire [temp_w*6-1:0] c1040ibus;
wire [data_w*6-1:0] c1040obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1040 ( .en(en), .clk(clk), .rst(rst), .q(c1040ibus), .r(c1040obus));
wire [temp_w*6-1:0] c1041ibus;
wire [data_w*6-1:0] c1041obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1041 ( .en(en), .clk(clk), .rst(rst), .q(c1041ibus), .r(c1041obus));
wire [temp_w*6-1:0] c1042ibus;
wire [data_w*6-1:0] c1042obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1042 ( .en(en), .clk(clk), .rst(rst), .q(c1042ibus), .r(c1042obus));
wire [temp_w*6-1:0] c1043ibus;
wire [data_w*6-1:0] c1043obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1043 ( .en(en), .clk(clk), .rst(rst), .q(c1043ibus), .r(c1043obus));
wire [temp_w*6-1:0] c1044ibus;
wire [data_w*6-1:0] c1044obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1044 ( .en(en), .clk(clk), .rst(rst), .q(c1044ibus), .r(c1044obus));
wire [temp_w*6-1:0] c1045ibus;
wire [data_w*6-1:0] c1045obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1045 ( .en(en), .clk(clk), .rst(rst), .q(c1045ibus), .r(c1045obus));
wire [temp_w*6-1:0] c1046ibus;
wire [data_w*6-1:0] c1046obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1046 ( .en(en), .clk(clk), .rst(rst), .q(c1046ibus), .r(c1046obus));
wire [temp_w*6-1:0] c1047ibus;
wire [data_w*6-1:0] c1047obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1047 ( .en(en), .clk(clk), .rst(rst), .q(c1047ibus), .r(c1047obus));
wire [temp_w*6-1:0] c1048ibus;
wire [data_w*6-1:0] c1048obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1048 ( .en(en), .clk(clk), .rst(rst), .q(c1048ibus), .r(c1048obus));
wire [temp_w*6-1:0] c1049ibus;
wire [data_w*6-1:0] c1049obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1049 ( .en(en), .clk(clk), .rst(rst), .q(c1049ibus), .r(c1049obus));
wire [temp_w*6-1:0] c1050ibus;
wire [data_w*6-1:0] c1050obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1050 ( .en(en), .clk(clk), .rst(rst), .q(c1050ibus), .r(c1050obus));
wire [temp_w*6-1:0] c1051ibus;
wire [data_w*6-1:0] c1051obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1051 ( .en(en), .clk(clk), .rst(rst), .q(c1051ibus), .r(c1051obus));
wire [temp_w*6-1:0] c1052ibus;
wire [data_w*6-1:0] c1052obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1052 ( .en(en), .clk(clk), .rst(rst), .q(c1052ibus), .r(c1052obus));
wire [temp_w*6-1:0] c1053ibus;
wire [data_w*6-1:0] c1053obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1053 ( .en(en), .clk(clk), .rst(rst), .q(c1053ibus), .r(c1053obus));
wire [temp_w*6-1:0] c1054ibus;
wire [data_w*6-1:0] c1054obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1054 ( .en(en), .clk(clk), .rst(rst), .q(c1054ibus), .r(c1054obus));
wire [temp_w*6-1:0] c1055ibus;
wire [data_w*6-1:0] c1055obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1055 ( .en(en), .clk(clk), .rst(rst), .q(c1055ibus), .r(c1055obus));
wire [temp_w*6-1:0] c1056ibus;
wire [data_w*6-1:0] c1056obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1056 ( .en(en), .clk(clk), .rst(rst), .q(c1056ibus), .r(c1056obus));
wire [temp_w*6-1:0] c1057ibus;
wire [data_w*6-1:0] c1057obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1057 ( .en(en), .clk(clk), .rst(rst), .q(c1057ibus), .r(c1057obus));
wire [temp_w*6-1:0] c1058ibus;
wire [data_w*6-1:0] c1058obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1058 ( .en(en), .clk(clk), .rst(rst), .q(c1058ibus), .r(c1058obus));
wire [temp_w*6-1:0] c1059ibus;
wire [data_w*6-1:0] c1059obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1059 ( .en(en), .clk(clk), .rst(rst), .q(c1059ibus), .r(c1059obus));
wire [temp_w*6-1:0] c1060ibus;
wire [data_w*6-1:0] c1060obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1060 ( .en(en), .clk(clk), .rst(rst), .q(c1060ibus), .r(c1060obus));
wire [temp_w*6-1:0] c1061ibus;
wire [data_w*6-1:0] c1061obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1061 ( .en(en), .clk(clk), .rst(rst), .q(c1061ibus), .r(c1061obus));
wire [temp_w*6-1:0] c1062ibus;
wire [data_w*6-1:0] c1062obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1062 ( .en(en), .clk(clk), .rst(rst), .q(c1062ibus), .r(c1062obus));
wire [temp_w*6-1:0] c1063ibus;
wire [data_w*6-1:0] c1063obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1063 ( .en(en), .clk(clk), .rst(rst), .q(c1063ibus), .r(c1063obus));
wire [temp_w*6-1:0] c1064ibus;
wire [data_w*6-1:0] c1064obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1064 ( .en(en), .clk(clk), .rst(rst), .q(c1064ibus), .r(c1064obus));
wire [temp_w*6-1:0] c1065ibus;
wire [data_w*6-1:0] c1065obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1065 ( .en(en), .clk(clk), .rst(rst), .q(c1065ibus), .r(c1065obus));
wire [temp_w*6-1:0] c1066ibus;
wire [data_w*6-1:0] c1066obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1066 ( .en(en), .clk(clk), .rst(rst), .q(c1066ibus), .r(c1066obus));
wire [temp_w*6-1:0] c1067ibus;
wire [data_w*6-1:0] c1067obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1067 ( .en(en), .clk(clk), .rst(rst), .q(c1067ibus), .r(c1067obus));
wire [temp_w*6-1:0] c1068ibus;
wire [data_w*6-1:0] c1068obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1068 ( .en(en), .clk(clk), .rst(rst), .q(c1068ibus), .r(c1068obus));
wire [temp_w*6-1:0] c1069ibus;
wire [data_w*6-1:0] c1069obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1069 ( .en(en), .clk(clk), .rst(rst), .q(c1069ibus), .r(c1069obus));
wire [temp_w*6-1:0] c1070ibus;
wire [data_w*6-1:0] c1070obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1070 ( .en(en), .clk(clk), .rst(rst), .q(c1070ibus), .r(c1070obus));
wire [temp_w*6-1:0] c1071ibus;
wire [data_w*6-1:0] c1071obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1071 ( .en(en), .clk(clk), .rst(rst), .q(c1071ibus), .r(c1071obus));
wire [temp_w*6-1:0] c1072ibus;
wire [data_w*6-1:0] c1072obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1072 ( .en(en), .clk(clk), .rst(rst), .q(c1072ibus), .r(c1072obus));
wire [temp_w*6-1:0] c1073ibus;
wire [data_w*6-1:0] c1073obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1073 ( .en(en), .clk(clk), .rst(rst), .q(c1073ibus), .r(c1073obus));
wire [temp_w*6-1:0] c1074ibus;
wire [data_w*6-1:0] c1074obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1074 ( .en(en), .clk(clk), .rst(rst), .q(c1074ibus), .r(c1074obus));
wire [temp_w*6-1:0] c1075ibus;
wire [data_w*6-1:0] c1075obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1075 ( .en(en), .clk(clk), .rst(rst), .q(c1075ibus), .r(c1075obus));
wire [temp_w*6-1:0] c1076ibus;
wire [data_w*6-1:0] c1076obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1076 ( .en(en), .clk(clk), .rst(rst), .q(c1076ibus), .r(c1076obus));
wire [temp_w*6-1:0] c1077ibus;
wire [data_w*6-1:0] c1077obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1077 ( .en(en), .clk(clk), .rst(rst), .q(c1077ibus), .r(c1077obus));
wire [temp_w*6-1:0] c1078ibus;
wire [data_w*6-1:0] c1078obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1078 ( .en(en), .clk(clk), .rst(rst), .q(c1078ibus), .r(c1078obus));
wire [temp_w*6-1:0] c1079ibus;
wire [data_w*6-1:0] c1079obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1079 ( .en(en), .clk(clk), .rst(rst), .q(c1079ibus), .r(c1079obus));
wire [temp_w*6-1:0] c1080ibus;
wire [data_w*6-1:0] c1080obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1080 ( .en(en), .clk(clk), .rst(rst), .q(c1080ibus), .r(c1080obus));
wire [temp_w*6-1:0] c1081ibus;
wire [data_w*6-1:0] c1081obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1081 ( .en(en), .clk(clk), .rst(rst), .q(c1081ibus), .r(c1081obus));
wire [temp_w*6-1:0] c1082ibus;
wire [data_w*6-1:0] c1082obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1082 ( .en(en), .clk(clk), .rst(rst), .q(c1082ibus), .r(c1082obus));
wire [temp_w*6-1:0] c1083ibus;
wire [data_w*6-1:0] c1083obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1083 ( .en(en), .clk(clk), .rst(rst), .q(c1083ibus), .r(c1083obus));
wire [temp_w*6-1:0] c1084ibus;
wire [data_w*6-1:0] c1084obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1084 ( .en(en), .clk(clk), .rst(rst), .q(c1084ibus), .r(c1084obus));
wire [temp_w*6-1:0] c1085ibus;
wire [data_w*6-1:0] c1085obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1085 ( .en(en), .clk(clk), .rst(rst), .q(c1085ibus), .r(c1085obus));
wire [temp_w*6-1:0] c1086ibus;
wire [data_w*6-1:0] c1086obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1086 ( .en(en), .clk(clk), .rst(rst), .q(c1086ibus), .r(c1086obus));
wire [temp_w*6-1:0] c1087ibus;
wire [data_w*6-1:0] c1087obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1087 ( .en(en), .clk(clk), .rst(rst), .q(c1087ibus), .r(c1087obus));
wire [temp_w*6-1:0] c1088ibus;
wire [data_w*6-1:0] c1088obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1088 ( .en(en), .clk(clk), .rst(rst), .q(c1088ibus), .r(c1088obus));
wire [temp_w*6-1:0] c1089ibus;
wire [data_w*6-1:0] c1089obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1089 ( .en(en), .clk(clk), .rst(rst), .q(c1089ibus), .r(c1089obus));
wire [temp_w*6-1:0] c1090ibus;
wire [data_w*6-1:0] c1090obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1090 ( .en(en), .clk(clk), .rst(rst), .q(c1090ibus), .r(c1090obus));
wire [temp_w*6-1:0] c1091ibus;
wire [data_w*6-1:0] c1091obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1091 ( .en(en), .clk(clk), .rst(rst), .q(c1091ibus), .r(c1091obus));
wire [temp_w*6-1:0] c1092ibus;
wire [data_w*6-1:0] c1092obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1092 ( .en(en), .clk(clk), .rst(rst), .q(c1092ibus), .r(c1092obus));
wire [temp_w*6-1:0] c1093ibus;
wire [data_w*6-1:0] c1093obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1093 ( .en(en), .clk(clk), .rst(rst), .q(c1093ibus), .r(c1093obus));
wire [temp_w*6-1:0] c1094ibus;
wire [data_w*6-1:0] c1094obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1094 ( .en(en), .clk(clk), .rst(rst), .q(c1094ibus), .r(c1094obus));
wire [temp_w*6-1:0] c1095ibus;
wire [data_w*6-1:0] c1095obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1095 ( .en(en), .clk(clk), .rst(rst), .q(c1095ibus), .r(c1095obus));
wire [temp_w*6-1:0] c1096ibus;
wire [data_w*6-1:0] c1096obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1096 ( .en(en), .clk(clk), .rst(rst), .q(c1096ibus), .r(c1096obus));
wire [temp_w*6-1:0] c1097ibus;
wire [data_w*6-1:0] c1097obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1097 ( .en(en), .clk(clk), .rst(rst), .q(c1097ibus), .r(c1097obus));
wire [temp_w*6-1:0] c1098ibus;
wire [data_w*6-1:0] c1098obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1098 ( .en(en), .clk(clk), .rst(rst), .q(c1098ibus), .r(c1098obus));
wire [temp_w*6-1:0] c1099ibus;
wire [data_w*6-1:0] c1099obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1099 ( .en(en), .clk(clk), .rst(rst), .q(c1099ibus), .r(c1099obus));
wire [temp_w*6-1:0] c1100ibus;
wire [data_w*6-1:0] c1100obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1100 ( .en(en), .clk(clk), .rst(rst), .q(c1100ibus), .r(c1100obus));
wire [temp_w*6-1:0] c1101ibus;
wire [data_w*6-1:0] c1101obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1101 ( .en(en), .clk(clk), .rst(rst), .q(c1101ibus), .r(c1101obus));
wire [temp_w*6-1:0] c1102ibus;
wire [data_w*6-1:0] c1102obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1102 ( .en(en), .clk(clk), .rst(rst), .q(c1102ibus), .r(c1102obus));
wire [temp_w*6-1:0] c1103ibus;
wire [data_w*6-1:0] c1103obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1103 ( .en(en), .clk(clk), .rst(rst), .q(c1103ibus), .r(c1103obus));
wire [temp_w*6-1:0] c1104ibus;
wire [data_w*6-1:0] c1104obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1104 ( .en(en), .clk(clk), .rst(rst), .q(c1104ibus), .r(c1104obus));
wire [temp_w*6-1:0] c1105ibus;
wire [data_w*6-1:0] c1105obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1105 ( .en(en), .clk(clk), .rst(rst), .q(c1105ibus), .r(c1105obus));
wire [temp_w*6-1:0] c1106ibus;
wire [data_w*6-1:0] c1106obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1106 ( .en(en), .clk(clk), .rst(rst), .q(c1106ibus), .r(c1106obus));
wire [temp_w*6-1:0] c1107ibus;
wire [data_w*6-1:0] c1107obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1107 ( .en(en), .clk(clk), .rst(rst), .q(c1107ibus), .r(c1107obus));
wire [temp_w*6-1:0] c1108ibus;
wire [data_w*6-1:0] c1108obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1108 ( .en(en), .clk(clk), .rst(rst), .q(c1108ibus), .r(c1108obus));
wire [temp_w*6-1:0] c1109ibus;
wire [data_w*6-1:0] c1109obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1109 ( .en(en), .clk(clk), .rst(rst), .q(c1109ibus), .r(c1109obus));
wire [temp_w*6-1:0] c1110ibus;
wire [data_w*6-1:0] c1110obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1110 ( .en(en), .clk(clk), .rst(rst), .q(c1110ibus), .r(c1110obus));
wire [temp_w*6-1:0] c1111ibus;
wire [data_w*6-1:0] c1111obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1111 ( .en(en), .clk(clk), .rst(rst), .q(c1111ibus), .r(c1111obus));
wire [temp_w*6-1:0] c1112ibus;
wire [data_w*6-1:0] c1112obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1112 ( .en(en), .clk(clk), .rst(rst), .q(c1112ibus), .r(c1112obus));
wire [temp_w*6-1:0] c1113ibus;
wire [data_w*6-1:0] c1113obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1113 ( .en(en), .clk(clk), .rst(rst), .q(c1113ibus), .r(c1113obus));
wire [temp_w*6-1:0] c1114ibus;
wire [data_w*6-1:0] c1114obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1114 ( .en(en), .clk(clk), .rst(rst), .q(c1114ibus), .r(c1114obus));
wire [temp_w*6-1:0] c1115ibus;
wire [data_w*6-1:0] c1115obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1115 ( .en(en), .clk(clk), .rst(rst), .q(c1115ibus), .r(c1115obus));
wire [temp_w*6-1:0] c1116ibus;
wire [data_w*6-1:0] c1116obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1116 ( .en(en), .clk(clk), .rst(rst), .q(c1116ibus), .r(c1116obus));
wire [temp_w*6-1:0] c1117ibus;
wire [data_w*6-1:0] c1117obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1117 ( .en(en), .clk(clk), .rst(rst), .q(c1117ibus), .r(c1117obus));
wire [temp_w*6-1:0] c1118ibus;
wire [data_w*6-1:0] c1118obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1118 ( .en(en), .clk(clk), .rst(rst), .q(c1118ibus), .r(c1118obus));
wire [temp_w*6-1:0] c1119ibus;
wire [data_w*6-1:0] c1119obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1119 ( .en(en), .clk(clk), .rst(rst), .q(c1119ibus), .r(c1119obus));
wire [temp_w*6-1:0] c1120ibus;
wire [data_w*6-1:0] c1120obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1120 ( .en(en), .clk(clk), .rst(rst), .q(c1120ibus), .r(c1120obus));
wire [temp_w*6-1:0] c1121ibus;
wire [data_w*6-1:0] c1121obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1121 ( .en(en), .clk(clk), .rst(rst), .q(c1121ibus), .r(c1121obus));
wire [temp_w*6-1:0] c1122ibus;
wire [data_w*6-1:0] c1122obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1122 ( .en(en), .clk(clk), .rst(rst), .q(c1122ibus), .r(c1122obus));
wire [temp_w*6-1:0] c1123ibus;
wire [data_w*6-1:0] c1123obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1123 ( .en(en), .clk(clk), .rst(rst), .q(c1123ibus), .r(c1123obus));
wire [temp_w*6-1:0] c1124ibus;
wire [data_w*6-1:0] c1124obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1124 ( .en(en), .clk(clk), .rst(rst), .q(c1124ibus), .r(c1124obus));
wire [temp_w*6-1:0] c1125ibus;
wire [data_w*6-1:0] c1125obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1125 ( .en(en), .clk(clk), .rst(rst), .q(c1125ibus), .r(c1125obus));
wire [temp_w*6-1:0] c1126ibus;
wire [data_w*6-1:0] c1126obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1126 ( .en(en), .clk(clk), .rst(rst), .q(c1126ibus), .r(c1126obus));
wire [temp_w*6-1:0] c1127ibus;
wire [data_w*6-1:0] c1127obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1127 ( .en(en), .clk(clk), .rst(rst), .q(c1127ibus), .r(c1127obus));
wire [temp_w*6-1:0] c1128ibus;
wire [data_w*6-1:0] c1128obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1128 ( .en(en), .clk(clk), .rst(rst), .q(c1128ibus), .r(c1128obus));
wire [temp_w*6-1:0] c1129ibus;
wire [data_w*6-1:0] c1129obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1129 ( .en(en), .clk(clk), .rst(rst), .q(c1129ibus), .r(c1129obus));
wire [temp_w*6-1:0] c1130ibus;
wire [data_w*6-1:0] c1130obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1130 ( .en(en), .clk(clk), .rst(rst), .q(c1130ibus), .r(c1130obus));
wire [temp_w*6-1:0] c1131ibus;
wire [data_w*6-1:0] c1131obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1131 ( .en(en), .clk(clk), .rst(rst), .q(c1131ibus), .r(c1131obus));
wire [temp_w*6-1:0] c1132ibus;
wire [data_w*6-1:0] c1132obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1132 ( .en(en), .clk(clk), .rst(rst), .q(c1132ibus), .r(c1132obus));
wire [temp_w*6-1:0] c1133ibus;
wire [data_w*6-1:0] c1133obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1133 ( .en(en), .clk(clk), .rst(rst), .q(c1133ibus), .r(c1133obus));
wire [temp_w*6-1:0] c1134ibus;
wire [data_w*6-1:0] c1134obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1134 ( .en(en), .clk(clk), .rst(rst), .q(c1134ibus), .r(c1134obus));
wire [temp_w*6-1:0] c1135ibus;
wire [data_w*6-1:0] c1135obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1135 ( .en(en), .clk(clk), .rst(rst), .q(c1135ibus), .r(c1135obus));
wire [temp_w*6-1:0] c1136ibus;
wire [data_w*6-1:0] c1136obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1136 ( .en(en), .clk(clk), .rst(rst), .q(c1136ibus), .r(c1136obus));
wire [temp_w*6-1:0] c1137ibus;
wire [data_w*6-1:0] c1137obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1137 ( .en(en), .clk(clk), .rst(rst), .q(c1137ibus), .r(c1137obus));
wire [temp_w*6-1:0] c1138ibus;
wire [data_w*6-1:0] c1138obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1138 ( .en(en), .clk(clk), .rst(rst), .q(c1138ibus), .r(c1138obus));
wire [temp_w*6-1:0] c1139ibus;
wire [data_w*6-1:0] c1139obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1139 ( .en(en), .clk(clk), .rst(rst), .q(c1139ibus), .r(c1139obus));
wire [temp_w*6-1:0] c1140ibus;
wire [data_w*6-1:0] c1140obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1140 ( .en(en), .clk(clk), .rst(rst), .q(c1140ibus), .r(c1140obus));
wire [temp_w*6-1:0] c1141ibus;
wire [data_w*6-1:0] c1141obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1141 ( .en(en), .clk(clk), .rst(rst), .q(c1141ibus), .r(c1141obus));
wire [temp_w*6-1:0] c1142ibus;
wire [data_w*6-1:0] c1142obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1142 ( .en(en), .clk(clk), .rst(rst), .q(c1142ibus), .r(c1142obus));
wire [temp_w*6-1:0] c1143ibus;
wire [data_w*6-1:0] c1143obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1143 ( .en(en), .clk(clk), .rst(rst), .q(c1143ibus), .r(c1143obus));
wire [temp_w*6-1:0] c1144ibus;
wire [data_w*6-1:0] c1144obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1144 ( .en(en), .clk(clk), .rst(rst), .q(c1144ibus), .r(c1144obus));
wire [temp_w*6-1:0] c1145ibus;
wire [data_w*6-1:0] c1145obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1145 ( .en(en), .clk(clk), .rst(rst), .q(c1145ibus), .r(c1145obus));
wire [temp_w*6-1:0] c1146ibus;
wire [data_w*6-1:0] c1146obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1146 ( .en(en), .clk(clk), .rst(rst), .q(c1146ibus), .r(c1146obus));
wire [temp_w*6-1:0] c1147ibus;
wire [data_w*6-1:0] c1147obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1147 ( .en(en), .clk(clk), .rst(rst), .q(c1147ibus), .r(c1147obus));
wire [temp_w*6-1:0] c1148ibus;
wire [data_w*6-1:0] c1148obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1148 ( .en(en), .clk(clk), .rst(rst), .q(c1148ibus), .r(c1148obus));
wire [temp_w*6-1:0] c1149ibus;
wire [data_w*6-1:0] c1149obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1149 ( .en(en), .clk(clk), .rst(rst), .q(c1149ibus), .r(c1149obus));
wire [temp_w*6-1:0] c1150ibus;
wire [data_w*6-1:0] c1150obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1150 ( .en(en), .clk(clk), .rst(rst), .q(c1150ibus), .r(c1150obus));
wire [temp_w*6-1:0] c1151ibus;
wire [data_w*6-1:0] c1151obus;
cnu #(.res_w(data_w), .ext_w(ext_w), .D(6), .idx_w(idx_w)) CNU1151 ( .en(en), .clk(clk), .rst(rst), .q(c1151ibus), .r(c1151obus));

wire [data_w*3-1:0] v0ibus;
wire [temp_w*3-1:0] v0obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU0 (.l(l[0*data_w +:data_w]), .r(v0ibus), .q(v0obus), .dec(dec[0]));
wire [data_w*3-1:0] v1ibus;
wire [temp_w*3-1:0] v1obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1 (.l(l[1*data_w +:data_w]), .r(v1ibus), .q(v1obus), .dec(dec[1]));
wire [data_w*3-1:0] v2ibus;
wire [temp_w*3-1:0] v2obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU2 (.l(l[2*data_w +:data_w]), .r(v2ibus), .q(v2obus), .dec(dec[2]));
wire [data_w*3-1:0] v3ibus;
wire [temp_w*3-1:0] v3obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU3 (.l(l[3*data_w +:data_w]), .r(v3ibus), .q(v3obus), .dec(dec[3]));
wire [data_w*3-1:0] v4ibus;
wire [temp_w*3-1:0] v4obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU4 (.l(l[4*data_w +:data_w]), .r(v4ibus), .q(v4obus), .dec(dec[4]));
wire [data_w*3-1:0] v5ibus;
wire [temp_w*3-1:0] v5obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU5 (.l(l[5*data_w +:data_w]), .r(v5ibus), .q(v5obus), .dec(dec[5]));
wire [data_w*3-1:0] v6ibus;
wire [temp_w*3-1:0] v6obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU6 (.l(l[6*data_w +:data_w]), .r(v6ibus), .q(v6obus), .dec(dec[6]));
wire [data_w*3-1:0] v7ibus;
wire [temp_w*3-1:0] v7obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU7 (.l(l[7*data_w +:data_w]), .r(v7ibus), .q(v7obus), .dec(dec[7]));
wire [data_w*3-1:0] v8ibus;
wire [temp_w*3-1:0] v8obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU8 (.l(l[8*data_w +:data_w]), .r(v8ibus), .q(v8obus), .dec(dec[8]));
wire [data_w*3-1:0] v9ibus;
wire [temp_w*3-1:0] v9obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU9 (.l(l[9*data_w +:data_w]), .r(v9ibus), .q(v9obus), .dec(dec[9]));
wire [data_w*3-1:0] v10ibus;
wire [temp_w*3-1:0] v10obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU10 (.l(l[10*data_w +:data_w]), .r(v10ibus), .q(v10obus), .dec(dec[10]));
wire [data_w*3-1:0] v11ibus;
wire [temp_w*3-1:0] v11obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU11 (.l(l[11*data_w +:data_w]), .r(v11ibus), .q(v11obus), .dec(dec[11]));
wire [data_w*3-1:0] v12ibus;
wire [temp_w*3-1:0] v12obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU12 (.l(l[12*data_w +:data_w]), .r(v12ibus), .q(v12obus), .dec(dec[12]));
wire [data_w*3-1:0] v13ibus;
wire [temp_w*3-1:0] v13obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU13 (.l(l[13*data_w +:data_w]), .r(v13ibus), .q(v13obus), .dec(dec[13]));
wire [data_w*3-1:0] v14ibus;
wire [temp_w*3-1:0] v14obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU14 (.l(l[14*data_w +:data_w]), .r(v14ibus), .q(v14obus), .dec(dec[14]));
wire [data_w*3-1:0] v15ibus;
wire [temp_w*3-1:0] v15obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU15 (.l(l[15*data_w +:data_w]), .r(v15ibus), .q(v15obus), .dec(dec[15]));
wire [data_w*3-1:0] v16ibus;
wire [temp_w*3-1:0] v16obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU16 (.l(l[16*data_w +:data_w]), .r(v16ibus), .q(v16obus), .dec(dec[16]));
wire [data_w*3-1:0] v17ibus;
wire [temp_w*3-1:0] v17obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU17 (.l(l[17*data_w +:data_w]), .r(v17ibus), .q(v17obus), .dec(dec[17]));
wire [data_w*3-1:0] v18ibus;
wire [temp_w*3-1:0] v18obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU18 (.l(l[18*data_w +:data_w]), .r(v18ibus), .q(v18obus), .dec(dec[18]));
wire [data_w*3-1:0] v19ibus;
wire [temp_w*3-1:0] v19obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU19 (.l(l[19*data_w +:data_w]), .r(v19ibus), .q(v19obus), .dec(dec[19]));
wire [data_w*3-1:0] v20ibus;
wire [temp_w*3-1:0] v20obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU20 (.l(l[20*data_w +:data_w]), .r(v20ibus), .q(v20obus), .dec(dec[20]));
wire [data_w*3-1:0] v21ibus;
wire [temp_w*3-1:0] v21obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU21 (.l(l[21*data_w +:data_w]), .r(v21ibus), .q(v21obus), .dec(dec[21]));
wire [data_w*3-1:0] v22ibus;
wire [temp_w*3-1:0] v22obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU22 (.l(l[22*data_w +:data_w]), .r(v22ibus), .q(v22obus), .dec(dec[22]));
wire [data_w*3-1:0] v23ibus;
wire [temp_w*3-1:0] v23obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU23 (.l(l[23*data_w +:data_w]), .r(v23ibus), .q(v23obus), .dec(dec[23]));
wire [data_w*3-1:0] v24ibus;
wire [temp_w*3-1:0] v24obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU24 (.l(l[24*data_w +:data_w]), .r(v24ibus), .q(v24obus), .dec(dec[24]));
wire [data_w*3-1:0] v25ibus;
wire [temp_w*3-1:0] v25obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU25 (.l(l[25*data_w +:data_w]), .r(v25ibus), .q(v25obus), .dec(dec[25]));
wire [data_w*3-1:0] v26ibus;
wire [temp_w*3-1:0] v26obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU26 (.l(l[26*data_w +:data_w]), .r(v26ibus), .q(v26obus), .dec(dec[26]));
wire [data_w*3-1:0] v27ibus;
wire [temp_w*3-1:0] v27obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU27 (.l(l[27*data_w +:data_w]), .r(v27ibus), .q(v27obus), .dec(dec[27]));
wire [data_w*3-1:0] v28ibus;
wire [temp_w*3-1:0] v28obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU28 (.l(l[28*data_w +:data_w]), .r(v28ibus), .q(v28obus), .dec(dec[28]));
wire [data_w*3-1:0] v29ibus;
wire [temp_w*3-1:0] v29obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU29 (.l(l[29*data_w +:data_w]), .r(v29ibus), .q(v29obus), .dec(dec[29]));
wire [data_w*3-1:0] v30ibus;
wire [temp_w*3-1:0] v30obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU30 (.l(l[30*data_w +:data_w]), .r(v30ibus), .q(v30obus), .dec(dec[30]));
wire [data_w*3-1:0] v31ibus;
wire [temp_w*3-1:0] v31obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU31 (.l(l[31*data_w +:data_w]), .r(v31ibus), .q(v31obus), .dec(dec[31]));
wire [data_w*3-1:0] v32ibus;
wire [temp_w*3-1:0] v32obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU32 (.l(l[32*data_w +:data_w]), .r(v32ibus), .q(v32obus), .dec(dec[32]));
wire [data_w*3-1:0] v33ibus;
wire [temp_w*3-1:0] v33obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU33 (.l(l[33*data_w +:data_w]), .r(v33ibus), .q(v33obus), .dec(dec[33]));
wire [data_w*3-1:0] v34ibus;
wire [temp_w*3-1:0] v34obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU34 (.l(l[34*data_w +:data_w]), .r(v34ibus), .q(v34obus), .dec(dec[34]));
wire [data_w*3-1:0] v35ibus;
wire [temp_w*3-1:0] v35obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU35 (.l(l[35*data_w +:data_w]), .r(v35ibus), .q(v35obus), .dec(dec[35]));
wire [data_w*3-1:0] v36ibus;
wire [temp_w*3-1:0] v36obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU36 (.l(l[36*data_w +:data_w]), .r(v36ibus), .q(v36obus), .dec(dec[36]));
wire [data_w*3-1:0] v37ibus;
wire [temp_w*3-1:0] v37obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU37 (.l(l[37*data_w +:data_w]), .r(v37ibus), .q(v37obus), .dec(dec[37]));
wire [data_w*3-1:0] v38ibus;
wire [temp_w*3-1:0] v38obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU38 (.l(l[38*data_w +:data_w]), .r(v38ibus), .q(v38obus), .dec(dec[38]));
wire [data_w*3-1:0] v39ibus;
wire [temp_w*3-1:0] v39obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU39 (.l(l[39*data_w +:data_w]), .r(v39ibus), .q(v39obus), .dec(dec[39]));
wire [data_w*3-1:0] v40ibus;
wire [temp_w*3-1:0] v40obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU40 (.l(l[40*data_w +:data_w]), .r(v40ibus), .q(v40obus), .dec(dec[40]));
wire [data_w*3-1:0] v41ibus;
wire [temp_w*3-1:0] v41obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU41 (.l(l[41*data_w +:data_w]), .r(v41ibus), .q(v41obus), .dec(dec[41]));
wire [data_w*3-1:0] v42ibus;
wire [temp_w*3-1:0] v42obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU42 (.l(l[42*data_w +:data_w]), .r(v42ibus), .q(v42obus), .dec(dec[42]));
wire [data_w*3-1:0] v43ibus;
wire [temp_w*3-1:0] v43obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU43 (.l(l[43*data_w +:data_w]), .r(v43ibus), .q(v43obus), .dec(dec[43]));
wire [data_w*3-1:0] v44ibus;
wire [temp_w*3-1:0] v44obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU44 (.l(l[44*data_w +:data_w]), .r(v44ibus), .q(v44obus), .dec(dec[44]));
wire [data_w*3-1:0] v45ibus;
wire [temp_w*3-1:0] v45obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU45 (.l(l[45*data_w +:data_w]), .r(v45ibus), .q(v45obus), .dec(dec[45]));
wire [data_w*3-1:0] v46ibus;
wire [temp_w*3-1:0] v46obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU46 (.l(l[46*data_w +:data_w]), .r(v46ibus), .q(v46obus), .dec(dec[46]));
wire [data_w*3-1:0] v47ibus;
wire [temp_w*3-1:0] v47obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU47 (.l(l[47*data_w +:data_w]), .r(v47ibus), .q(v47obus), .dec(dec[47]));
wire [data_w*3-1:0] v48ibus;
wire [temp_w*3-1:0] v48obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU48 (.l(l[48*data_w +:data_w]), .r(v48ibus), .q(v48obus), .dec(dec[48]));
wire [data_w*3-1:0] v49ibus;
wire [temp_w*3-1:0] v49obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU49 (.l(l[49*data_w +:data_w]), .r(v49ibus), .q(v49obus), .dec(dec[49]));
wire [data_w*3-1:0] v50ibus;
wire [temp_w*3-1:0] v50obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU50 (.l(l[50*data_w +:data_w]), .r(v50ibus), .q(v50obus), .dec(dec[50]));
wire [data_w*3-1:0] v51ibus;
wire [temp_w*3-1:0] v51obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU51 (.l(l[51*data_w +:data_w]), .r(v51ibus), .q(v51obus), .dec(dec[51]));
wire [data_w*3-1:0] v52ibus;
wire [temp_w*3-1:0] v52obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU52 (.l(l[52*data_w +:data_w]), .r(v52ibus), .q(v52obus), .dec(dec[52]));
wire [data_w*3-1:0] v53ibus;
wire [temp_w*3-1:0] v53obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU53 (.l(l[53*data_w +:data_w]), .r(v53ibus), .q(v53obus), .dec(dec[53]));
wire [data_w*3-1:0] v54ibus;
wire [temp_w*3-1:0] v54obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU54 (.l(l[54*data_w +:data_w]), .r(v54ibus), .q(v54obus), .dec(dec[54]));
wire [data_w*3-1:0] v55ibus;
wire [temp_w*3-1:0] v55obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU55 (.l(l[55*data_w +:data_w]), .r(v55ibus), .q(v55obus), .dec(dec[55]));
wire [data_w*3-1:0] v56ibus;
wire [temp_w*3-1:0] v56obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU56 (.l(l[56*data_w +:data_w]), .r(v56ibus), .q(v56obus), .dec(dec[56]));
wire [data_w*3-1:0] v57ibus;
wire [temp_w*3-1:0] v57obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU57 (.l(l[57*data_w +:data_w]), .r(v57ibus), .q(v57obus), .dec(dec[57]));
wire [data_w*3-1:0] v58ibus;
wire [temp_w*3-1:0] v58obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU58 (.l(l[58*data_w +:data_w]), .r(v58ibus), .q(v58obus), .dec(dec[58]));
wire [data_w*3-1:0] v59ibus;
wire [temp_w*3-1:0] v59obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU59 (.l(l[59*data_w +:data_w]), .r(v59ibus), .q(v59obus), .dec(dec[59]));
wire [data_w*3-1:0] v60ibus;
wire [temp_w*3-1:0] v60obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU60 (.l(l[60*data_w +:data_w]), .r(v60ibus), .q(v60obus), .dec(dec[60]));
wire [data_w*3-1:0] v61ibus;
wire [temp_w*3-1:0] v61obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU61 (.l(l[61*data_w +:data_w]), .r(v61ibus), .q(v61obus), .dec(dec[61]));
wire [data_w*3-1:0] v62ibus;
wire [temp_w*3-1:0] v62obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU62 (.l(l[62*data_w +:data_w]), .r(v62ibus), .q(v62obus), .dec(dec[62]));
wire [data_w*3-1:0] v63ibus;
wire [temp_w*3-1:0] v63obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU63 (.l(l[63*data_w +:data_w]), .r(v63ibus), .q(v63obus), .dec(dec[63]));
wire [data_w*3-1:0] v64ibus;
wire [temp_w*3-1:0] v64obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU64 (.l(l[64*data_w +:data_w]), .r(v64ibus), .q(v64obus), .dec(dec[64]));
wire [data_w*3-1:0] v65ibus;
wire [temp_w*3-1:0] v65obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU65 (.l(l[65*data_w +:data_w]), .r(v65ibus), .q(v65obus), .dec(dec[65]));
wire [data_w*3-1:0] v66ibus;
wire [temp_w*3-1:0] v66obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU66 (.l(l[66*data_w +:data_w]), .r(v66ibus), .q(v66obus), .dec(dec[66]));
wire [data_w*3-1:0] v67ibus;
wire [temp_w*3-1:0] v67obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU67 (.l(l[67*data_w +:data_w]), .r(v67ibus), .q(v67obus), .dec(dec[67]));
wire [data_w*3-1:0] v68ibus;
wire [temp_w*3-1:0] v68obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU68 (.l(l[68*data_w +:data_w]), .r(v68ibus), .q(v68obus), .dec(dec[68]));
wire [data_w*3-1:0] v69ibus;
wire [temp_w*3-1:0] v69obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU69 (.l(l[69*data_w +:data_w]), .r(v69ibus), .q(v69obus), .dec(dec[69]));
wire [data_w*3-1:0] v70ibus;
wire [temp_w*3-1:0] v70obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU70 (.l(l[70*data_w +:data_w]), .r(v70ibus), .q(v70obus), .dec(dec[70]));
wire [data_w*3-1:0] v71ibus;
wire [temp_w*3-1:0] v71obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU71 (.l(l[71*data_w +:data_w]), .r(v71ibus), .q(v71obus), .dec(dec[71]));
wire [data_w*3-1:0] v72ibus;
wire [temp_w*3-1:0] v72obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU72 (.l(l[72*data_w +:data_w]), .r(v72ibus), .q(v72obus), .dec(dec[72]));
wire [data_w*3-1:0] v73ibus;
wire [temp_w*3-1:0] v73obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU73 (.l(l[73*data_w +:data_w]), .r(v73ibus), .q(v73obus), .dec(dec[73]));
wire [data_w*3-1:0] v74ibus;
wire [temp_w*3-1:0] v74obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU74 (.l(l[74*data_w +:data_w]), .r(v74ibus), .q(v74obus), .dec(dec[74]));
wire [data_w*3-1:0] v75ibus;
wire [temp_w*3-1:0] v75obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU75 (.l(l[75*data_w +:data_w]), .r(v75ibus), .q(v75obus), .dec(dec[75]));
wire [data_w*3-1:0] v76ibus;
wire [temp_w*3-1:0] v76obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU76 (.l(l[76*data_w +:data_w]), .r(v76ibus), .q(v76obus), .dec(dec[76]));
wire [data_w*3-1:0] v77ibus;
wire [temp_w*3-1:0] v77obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU77 (.l(l[77*data_w +:data_w]), .r(v77ibus), .q(v77obus), .dec(dec[77]));
wire [data_w*3-1:0] v78ibus;
wire [temp_w*3-1:0] v78obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU78 (.l(l[78*data_w +:data_w]), .r(v78ibus), .q(v78obus), .dec(dec[78]));
wire [data_w*3-1:0] v79ibus;
wire [temp_w*3-1:0] v79obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU79 (.l(l[79*data_w +:data_w]), .r(v79ibus), .q(v79obus), .dec(dec[79]));
wire [data_w*3-1:0] v80ibus;
wire [temp_w*3-1:0] v80obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU80 (.l(l[80*data_w +:data_w]), .r(v80ibus), .q(v80obus), .dec(dec[80]));
wire [data_w*3-1:0] v81ibus;
wire [temp_w*3-1:0] v81obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU81 (.l(l[81*data_w +:data_w]), .r(v81ibus), .q(v81obus), .dec(dec[81]));
wire [data_w*3-1:0] v82ibus;
wire [temp_w*3-1:0] v82obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU82 (.l(l[82*data_w +:data_w]), .r(v82ibus), .q(v82obus), .dec(dec[82]));
wire [data_w*3-1:0] v83ibus;
wire [temp_w*3-1:0] v83obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU83 (.l(l[83*data_w +:data_w]), .r(v83ibus), .q(v83obus), .dec(dec[83]));
wire [data_w*3-1:0] v84ibus;
wire [temp_w*3-1:0] v84obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU84 (.l(l[84*data_w +:data_w]), .r(v84ibus), .q(v84obus), .dec(dec[84]));
wire [data_w*3-1:0] v85ibus;
wire [temp_w*3-1:0] v85obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU85 (.l(l[85*data_w +:data_w]), .r(v85ibus), .q(v85obus), .dec(dec[85]));
wire [data_w*3-1:0] v86ibus;
wire [temp_w*3-1:0] v86obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU86 (.l(l[86*data_w +:data_w]), .r(v86ibus), .q(v86obus), .dec(dec[86]));
wire [data_w*3-1:0] v87ibus;
wire [temp_w*3-1:0] v87obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU87 (.l(l[87*data_w +:data_w]), .r(v87ibus), .q(v87obus), .dec(dec[87]));
wire [data_w*3-1:0] v88ibus;
wire [temp_w*3-1:0] v88obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU88 (.l(l[88*data_w +:data_w]), .r(v88ibus), .q(v88obus), .dec(dec[88]));
wire [data_w*3-1:0] v89ibus;
wire [temp_w*3-1:0] v89obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU89 (.l(l[89*data_w +:data_w]), .r(v89ibus), .q(v89obus), .dec(dec[89]));
wire [data_w*3-1:0] v90ibus;
wire [temp_w*3-1:0] v90obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU90 (.l(l[90*data_w +:data_w]), .r(v90ibus), .q(v90obus), .dec(dec[90]));
wire [data_w*3-1:0] v91ibus;
wire [temp_w*3-1:0] v91obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU91 (.l(l[91*data_w +:data_w]), .r(v91ibus), .q(v91obus), .dec(dec[91]));
wire [data_w*3-1:0] v92ibus;
wire [temp_w*3-1:0] v92obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU92 (.l(l[92*data_w +:data_w]), .r(v92ibus), .q(v92obus), .dec(dec[92]));
wire [data_w*3-1:0] v93ibus;
wire [temp_w*3-1:0] v93obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU93 (.l(l[93*data_w +:data_w]), .r(v93ibus), .q(v93obus), .dec(dec[93]));
wire [data_w*3-1:0] v94ibus;
wire [temp_w*3-1:0] v94obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU94 (.l(l[94*data_w +:data_w]), .r(v94ibus), .q(v94obus), .dec(dec[94]));
wire [data_w*3-1:0] v95ibus;
wire [temp_w*3-1:0] v95obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU95 (.l(l[95*data_w +:data_w]), .r(v95ibus), .q(v95obus), .dec(dec[95]));
wire [data_w*3-1:0] v96ibus;
wire [temp_w*3-1:0] v96obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU96 (.l(l[96*data_w +:data_w]), .r(v96ibus), .q(v96obus), .dec(dec[96]));
wire [data_w*3-1:0] v97ibus;
wire [temp_w*3-1:0] v97obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU97 (.l(l[97*data_w +:data_w]), .r(v97ibus), .q(v97obus), .dec(dec[97]));
wire [data_w*3-1:0] v98ibus;
wire [temp_w*3-1:0] v98obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU98 (.l(l[98*data_w +:data_w]), .r(v98ibus), .q(v98obus), .dec(dec[98]));
wire [data_w*3-1:0] v99ibus;
wire [temp_w*3-1:0] v99obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU99 (.l(l[99*data_w +:data_w]), .r(v99ibus), .q(v99obus), .dec(dec[99]));
wire [data_w*3-1:0] v100ibus;
wire [temp_w*3-1:0] v100obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU100 (.l(l[100*data_w +:data_w]), .r(v100ibus), .q(v100obus), .dec(dec[100]));
wire [data_w*3-1:0] v101ibus;
wire [temp_w*3-1:0] v101obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU101 (.l(l[101*data_w +:data_w]), .r(v101ibus), .q(v101obus), .dec(dec[101]));
wire [data_w*3-1:0] v102ibus;
wire [temp_w*3-1:0] v102obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU102 (.l(l[102*data_w +:data_w]), .r(v102ibus), .q(v102obus), .dec(dec[102]));
wire [data_w*3-1:0] v103ibus;
wire [temp_w*3-1:0] v103obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU103 (.l(l[103*data_w +:data_w]), .r(v103ibus), .q(v103obus), .dec(dec[103]));
wire [data_w*3-1:0] v104ibus;
wire [temp_w*3-1:0] v104obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU104 (.l(l[104*data_w +:data_w]), .r(v104ibus), .q(v104obus), .dec(dec[104]));
wire [data_w*3-1:0] v105ibus;
wire [temp_w*3-1:0] v105obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU105 (.l(l[105*data_w +:data_w]), .r(v105ibus), .q(v105obus), .dec(dec[105]));
wire [data_w*3-1:0] v106ibus;
wire [temp_w*3-1:0] v106obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU106 (.l(l[106*data_w +:data_w]), .r(v106ibus), .q(v106obus), .dec(dec[106]));
wire [data_w*3-1:0] v107ibus;
wire [temp_w*3-1:0] v107obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU107 (.l(l[107*data_w +:data_w]), .r(v107ibus), .q(v107obus), .dec(dec[107]));
wire [data_w*3-1:0] v108ibus;
wire [temp_w*3-1:0] v108obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU108 (.l(l[108*data_w +:data_w]), .r(v108ibus), .q(v108obus), .dec(dec[108]));
wire [data_w*3-1:0] v109ibus;
wire [temp_w*3-1:0] v109obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU109 (.l(l[109*data_w +:data_w]), .r(v109ibus), .q(v109obus), .dec(dec[109]));
wire [data_w*3-1:0] v110ibus;
wire [temp_w*3-1:0] v110obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU110 (.l(l[110*data_w +:data_w]), .r(v110ibus), .q(v110obus), .dec(dec[110]));
wire [data_w*3-1:0] v111ibus;
wire [temp_w*3-1:0] v111obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU111 (.l(l[111*data_w +:data_w]), .r(v111ibus), .q(v111obus), .dec(dec[111]));
wire [data_w*3-1:0] v112ibus;
wire [temp_w*3-1:0] v112obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU112 (.l(l[112*data_w +:data_w]), .r(v112ibus), .q(v112obus), .dec(dec[112]));
wire [data_w*3-1:0] v113ibus;
wire [temp_w*3-1:0] v113obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU113 (.l(l[113*data_w +:data_w]), .r(v113ibus), .q(v113obus), .dec(dec[113]));
wire [data_w*3-1:0] v114ibus;
wire [temp_w*3-1:0] v114obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU114 (.l(l[114*data_w +:data_w]), .r(v114ibus), .q(v114obus), .dec(dec[114]));
wire [data_w*3-1:0] v115ibus;
wire [temp_w*3-1:0] v115obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU115 (.l(l[115*data_w +:data_w]), .r(v115ibus), .q(v115obus), .dec(dec[115]));
wire [data_w*3-1:0] v116ibus;
wire [temp_w*3-1:0] v116obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU116 (.l(l[116*data_w +:data_w]), .r(v116ibus), .q(v116obus), .dec(dec[116]));
wire [data_w*3-1:0] v117ibus;
wire [temp_w*3-1:0] v117obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU117 (.l(l[117*data_w +:data_w]), .r(v117ibus), .q(v117obus), .dec(dec[117]));
wire [data_w*3-1:0] v118ibus;
wire [temp_w*3-1:0] v118obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU118 (.l(l[118*data_w +:data_w]), .r(v118ibus), .q(v118obus), .dec(dec[118]));
wire [data_w*3-1:0] v119ibus;
wire [temp_w*3-1:0] v119obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU119 (.l(l[119*data_w +:data_w]), .r(v119ibus), .q(v119obus), .dec(dec[119]));
wire [data_w*3-1:0] v120ibus;
wire [temp_w*3-1:0] v120obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU120 (.l(l[120*data_w +:data_w]), .r(v120ibus), .q(v120obus), .dec(dec[120]));
wire [data_w*3-1:0] v121ibus;
wire [temp_w*3-1:0] v121obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU121 (.l(l[121*data_w +:data_w]), .r(v121ibus), .q(v121obus), .dec(dec[121]));
wire [data_w*3-1:0] v122ibus;
wire [temp_w*3-1:0] v122obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU122 (.l(l[122*data_w +:data_w]), .r(v122ibus), .q(v122obus), .dec(dec[122]));
wire [data_w*3-1:0] v123ibus;
wire [temp_w*3-1:0] v123obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU123 (.l(l[123*data_w +:data_w]), .r(v123ibus), .q(v123obus), .dec(dec[123]));
wire [data_w*3-1:0] v124ibus;
wire [temp_w*3-1:0] v124obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU124 (.l(l[124*data_w +:data_w]), .r(v124ibus), .q(v124obus), .dec(dec[124]));
wire [data_w*3-1:0] v125ibus;
wire [temp_w*3-1:0] v125obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU125 (.l(l[125*data_w +:data_w]), .r(v125ibus), .q(v125obus), .dec(dec[125]));
wire [data_w*3-1:0] v126ibus;
wire [temp_w*3-1:0] v126obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU126 (.l(l[126*data_w +:data_w]), .r(v126ibus), .q(v126obus), .dec(dec[126]));
wire [data_w*3-1:0] v127ibus;
wire [temp_w*3-1:0] v127obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU127 (.l(l[127*data_w +:data_w]), .r(v127ibus), .q(v127obus), .dec(dec[127]));
wire [data_w*3-1:0] v128ibus;
wire [temp_w*3-1:0] v128obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU128 (.l(l[128*data_w +:data_w]), .r(v128ibus), .q(v128obus), .dec(dec[128]));
wire [data_w*3-1:0] v129ibus;
wire [temp_w*3-1:0] v129obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU129 (.l(l[129*data_w +:data_w]), .r(v129ibus), .q(v129obus), .dec(dec[129]));
wire [data_w*3-1:0] v130ibus;
wire [temp_w*3-1:0] v130obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU130 (.l(l[130*data_w +:data_w]), .r(v130ibus), .q(v130obus), .dec(dec[130]));
wire [data_w*3-1:0] v131ibus;
wire [temp_w*3-1:0] v131obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU131 (.l(l[131*data_w +:data_w]), .r(v131ibus), .q(v131obus), .dec(dec[131]));
wire [data_w*3-1:0] v132ibus;
wire [temp_w*3-1:0] v132obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU132 (.l(l[132*data_w +:data_w]), .r(v132ibus), .q(v132obus), .dec(dec[132]));
wire [data_w*3-1:0] v133ibus;
wire [temp_w*3-1:0] v133obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU133 (.l(l[133*data_w +:data_w]), .r(v133ibus), .q(v133obus), .dec(dec[133]));
wire [data_w*3-1:0] v134ibus;
wire [temp_w*3-1:0] v134obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU134 (.l(l[134*data_w +:data_w]), .r(v134ibus), .q(v134obus), .dec(dec[134]));
wire [data_w*3-1:0] v135ibus;
wire [temp_w*3-1:0] v135obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU135 (.l(l[135*data_w +:data_w]), .r(v135ibus), .q(v135obus), .dec(dec[135]));
wire [data_w*3-1:0] v136ibus;
wire [temp_w*3-1:0] v136obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU136 (.l(l[136*data_w +:data_w]), .r(v136ibus), .q(v136obus), .dec(dec[136]));
wire [data_w*3-1:0] v137ibus;
wire [temp_w*3-1:0] v137obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU137 (.l(l[137*data_w +:data_w]), .r(v137ibus), .q(v137obus), .dec(dec[137]));
wire [data_w*3-1:0] v138ibus;
wire [temp_w*3-1:0] v138obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU138 (.l(l[138*data_w +:data_w]), .r(v138ibus), .q(v138obus), .dec(dec[138]));
wire [data_w*3-1:0] v139ibus;
wire [temp_w*3-1:0] v139obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU139 (.l(l[139*data_w +:data_w]), .r(v139ibus), .q(v139obus), .dec(dec[139]));
wire [data_w*3-1:0] v140ibus;
wire [temp_w*3-1:0] v140obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU140 (.l(l[140*data_w +:data_w]), .r(v140ibus), .q(v140obus), .dec(dec[140]));
wire [data_w*3-1:0] v141ibus;
wire [temp_w*3-1:0] v141obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU141 (.l(l[141*data_w +:data_w]), .r(v141ibus), .q(v141obus), .dec(dec[141]));
wire [data_w*3-1:0] v142ibus;
wire [temp_w*3-1:0] v142obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU142 (.l(l[142*data_w +:data_w]), .r(v142ibus), .q(v142obus), .dec(dec[142]));
wire [data_w*3-1:0] v143ibus;
wire [temp_w*3-1:0] v143obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU143 (.l(l[143*data_w +:data_w]), .r(v143ibus), .q(v143obus), .dec(dec[143]));
wire [data_w*3-1:0] v144ibus;
wire [temp_w*3-1:0] v144obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU144 (.l(l[144*data_w +:data_w]), .r(v144ibus), .q(v144obus), .dec(dec[144]));
wire [data_w*3-1:0] v145ibus;
wire [temp_w*3-1:0] v145obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU145 (.l(l[145*data_w +:data_w]), .r(v145ibus), .q(v145obus), .dec(dec[145]));
wire [data_w*3-1:0] v146ibus;
wire [temp_w*3-1:0] v146obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU146 (.l(l[146*data_w +:data_w]), .r(v146ibus), .q(v146obus), .dec(dec[146]));
wire [data_w*3-1:0] v147ibus;
wire [temp_w*3-1:0] v147obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU147 (.l(l[147*data_w +:data_w]), .r(v147ibus), .q(v147obus), .dec(dec[147]));
wire [data_w*3-1:0] v148ibus;
wire [temp_w*3-1:0] v148obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU148 (.l(l[148*data_w +:data_w]), .r(v148ibus), .q(v148obus), .dec(dec[148]));
wire [data_w*3-1:0] v149ibus;
wire [temp_w*3-1:0] v149obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU149 (.l(l[149*data_w +:data_w]), .r(v149ibus), .q(v149obus), .dec(dec[149]));
wire [data_w*3-1:0] v150ibus;
wire [temp_w*3-1:0] v150obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU150 (.l(l[150*data_w +:data_w]), .r(v150ibus), .q(v150obus), .dec(dec[150]));
wire [data_w*3-1:0] v151ibus;
wire [temp_w*3-1:0] v151obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU151 (.l(l[151*data_w +:data_w]), .r(v151ibus), .q(v151obus), .dec(dec[151]));
wire [data_w*3-1:0] v152ibus;
wire [temp_w*3-1:0] v152obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU152 (.l(l[152*data_w +:data_w]), .r(v152ibus), .q(v152obus), .dec(dec[152]));
wire [data_w*3-1:0] v153ibus;
wire [temp_w*3-1:0] v153obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU153 (.l(l[153*data_w +:data_w]), .r(v153ibus), .q(v153obus), .dec(dec[153]));
wire [data_w*3-1:0] v154ibus;
wire [temp_w*3-1:0] v154obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU154 (.l(l[154*data_w +:data_w]), .r(v154ibus), .q(v154obus), .dec(dec[154]));
wire [data_w*3-1:0] v155ibus;
wire [temp_w*3-1:0] v155obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU155 (.l(l[155*data_w +:data_w]), .r(v155ibus), .q(v155obus), .dec(dec[155]));
wire [data_w*3-1:0] v156ibus;
wire [temp_w*3-1:0] v156obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU156 (.l(l[156*data_w +:data_w]), .r(v156ibus), .q(v156obus), .dec(dec[156]));
wire [data_w*3-1:0] v157ibus;
wire [temp_w*3-1:0] v157obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU157 (.l(l[157*data_w +:data_w]), .r(v157ibus), .q(v157obus), .dec(dec[157]));
wire [data_w*3-1:0] v158ibus;
wire [temp_w*3-1:0] v158obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU158 (.l(l[158*data_w +:data_w]), .r(v158ibus), .q(v158obus), .dec(dec[158]));
wire [data_w*3-1:0] v159ibus;
wire [temp_w*3-1:0] v159obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU159 (.l(l[159*data_w +:data_w]), .r(v159ibus), .q(v159obus), .dec(dec[159]));
wire [data_w*3-1:0] v160ibus;
wire [temp_w*3-1:0] v160obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU160 (.l(l[160*data_w +:data_w]), .r(v160ibus), .q(v160obus), .dec(dec[160]));
wire [data_w*3-1:0] v161ibus;
wire [temp_w*3-1:0] v161obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU161 (.l(l[161*data_w +:data_w]), .r(v161ibus), .q(v161obus), .dec(dec[161]));
wire [data_w*3-1:0] v162ibus;
wire [temp_w*3-1:0] v162obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU162 (.l(l[162*data_w +:data_w]), .r(v162ibus), .q(v162obus), .dec(dec[162]));
wire [data_w*3-1:0] v163ibus;
wire [temp_w*3-1:0] v163obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU163 (.l(l[163*data_w +:data_w]), .r(v163ibus), .q(v163obus), .dec(dec[163]));
wire [data_w*3-1:0] v164ibus;
wire [temp_w*3-1:0] v164obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU164 (.l(l[164*data_w +:data_w]), .r(v164ibus), .q(v164obus), .dec(dec[164]));
wire [data_w*3-1:0] v165ibus;
wire [temp_w*3-1:0] v165obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU165 (.l(l[165*data_w +:data_w]), .r(v165ibus), .q(v165obus), .dec(dec[165]));
wire [data_w*3-1:0] v166ibus;
wire [temp_w*3-1:0] v166obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU166 (.l(l[166*data_w +:data_w]), .r(v166ibus), .q(v166obus), .dec(dec[166]));
wire [data_w*3-1:0] v167ibus;
wire [temp_w*3-1:0] v167obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU167 (.l(l[167*data_w +:data_w]), .r(v167ibus), .q(v167obus), .dec(dec[167]));
wire [data_w*3-1:0] v168ibus;
wire [temp_w*3-1:0] v168obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU168 (.l(l[168*data_w +:data_w]), .r(v168ibus), .q(v168obus), .dec(dec[168]));
wire [data_w*3-1:0] v169ibus;
wire [temp_w*3-1:0] v169obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU169 (.l(l[169*data_w +:data_w]), .r(v169ibus), .q(v169obus), .dec(dec[169]));
wire [data_w*3-1:0] v170ibus;
wire [temp_w*3-1:0] v170obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU170 (.l(l[170*data_w +:data_w]), .r(v170ibus), .q(v170obus), .dec(dec[170]));
wire [data_w*3-1:0] v171ibus;
wire [temp_w*3-1:0] v171obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU171 (.l(l[171*data_w +:data_w]), .r(v171ibus), .q(v171obus), .dec(dec[171]));
wire [data_w*3-1:0] v172ibus;
wire [temp_w*3-1:0] v172obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU172 (.l(l[172*data_w +:data_w]), .r(v172ibus), .q(v172obus), .dec(dec[172]));
wire [data_w*3-1:0] v173ibus;
wire [temp_w*3-1:0] v173obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU173 (.l(l[173*data_w +:data_w]), .r(v173ibus), .q(v173obus), .dec(dec[173]));
wire [data_w*3-1:0] v174ibus;
wire [temp_w*3-1:0] v174obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU174 (.l(l[174*data_w +:data_w]), .r(v174ibus), .q(v174obus), .dec(dec[174]));
wire [data_w*3-1:0] v175ibus;
wire [temp_w*3-1:0] v175obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU175 (.l(l[175*data_w +:data_w]), .r(v175ibus), .q(v175obus), .dec(dec[175]));
wire [data_w*3-1:0] v176ibus;
wire [temp_w*3-1:0] v176obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU176 (.l(l[176*data_w +:data_w]), .r(v176ibus), .q(v176obus), .dec(dec[176]));
wire [data_w*3-1:0] v177ibus;
wire [temp_w*3-1:0] v177obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU177 (.l(l[177*data_w +:data_w]), .r(v177ibus), .q(v177obus), .dec(dec[177]));
wire [data_w*3-1:0] v178ibus;
wire [temp_w*3-1:0] v178obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU178 (.l(l[178*data_w +:data_w]), .r(v178ibus), .q(v178obus), .dec(dec[178]));
wire [data_w*3-1:0] v179ibus;
wire [temp_w*3-1:0] v179obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU179 (.l(l[179*data_w +:data_w]), .r(v179ibus), .q(v179obus), .dec(dec[179]));
wire [data_w*3-1:0] v180ibus;
wire [temp_w*3-1:0] v180obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU180 (.l(l[180*data_w +:data_w]), .r(v180ibus), .q(v180obus), .dec(dec[180]));
wire [data_w*3-1:0] v181ibus;
wire [temp_w*3-1:0] v181obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU181 (.l(l[181*data_w +:data_w]), .r(v181ibus), .q(v181obus), .dec(dec[181]));
wire [data_w*3-1:0] v182ibus;
wire [temp_w*3-1:0] v182obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU182 (.l(l[182*data_w +:data_w]), .r(v182ibus), .q(v182obus), .dec(dec[182]));
wire [data_w*3-1:0] v183ibus;
wire [temp_w*3-1:0] v183obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU183 (.l(l[183*data_w +:data_w]), .r(v183ibus), .q(v183obus), .dec(dec[183]));
wire [data_w*3-1:0] v184ibus;
wire [temp_w*3-1:0] v184obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU184 (.l(l[184*data_w +:data_w]), .r(v184ibus), .q(v184obus), .dec(dec[184]));
wire [data_w*3-1:0] v185ibus;
wire [temp_w*3-1:0] v185obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU185 (.l(l[185*data_w +:data_w]), .r(v185ibus), .q(v185obus), .dec(dec[185]));
wire [data_w*3-1:0] v186ibus;
wire [temp_w*3-1:0] v186obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU186 (.l(l[186*data_w +:data_w]), .r(v186ibus), .q(v186obus), .dec(dec[186]));
wire [data_w*3-1:0] v187ibus;
wire [temp_w*3-1:0] v187obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU187 (.l(l[187*data_w +:data_w]), .r(v187ibus), .q(v187obus), .dec(dec[187]));
wire [data_w*3-1:0] v188ibus;
wire [temp_w*3-1:0] v188obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU188 (.l(l[188*data_w +:data_w]), .r(v188ibus), .q(v188obus), .dec(dec[188]));
wire [data_w*3-1:0] v189ibus;
wire [temp_w*3-1:0] v189obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU189 (.l(l[189*data_w +:data_w]), .r(v189ibus), .q(v189obus), .dec(dec[189]));
wire [data_w*3-1:0] v190ibus;
wire [temp_w*3-1:0] v190obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU190 (.l(l[190*data_w +:data_w]), .r(v190ibus), .q(v190obus), .dec(dec[190]));
wire [data_w*3-1:0] v191ibus;
wire [temp_w*3-1:0] v191obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU191 (.l(l[191*data_w +:data_w]), .r(v191ibus), .q(v191obus), .dec(dec[191]));
wire [data_w*6-1:0] v192ibus;
wire [temp_w*6-1:0] v192obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU192 (.l(l[192*data_w +:data_w]), .r(v192ibus), .q(v192obus), .dec(dec[192]));
wire [data_w*6-1:0] v193ibus;
wire [temp_w*6-1:0] v193obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU193 (.l(l[193*data_w +:data_w]), .r(v193ibus), .q(v193obus), .dec(dec[193]));
wire [data_w*6-1:0] v194ibus;
wire [temp_w*6-1:0] v194obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU194 (.l(l[194*data_w +:data_w]), .r(v194ibus), .q(v194obus), .dec(dec[194]));
wire [data_w*6-1:0] v195ibus;
wire [temp_w*6-1:0] v195obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU195 (.l(l[195*data_w +:data_w]), .r(v195ibus), .q(v195obus), .dec(dec[195]));
wire [data_w*6-1:0] v196ibus;
wire [temp_w*6-1:0] v196obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU196 (.l(l[196*data_w +:data_w]), .r(v196ibus), .q(v196obus), .dec(dec[196]));
wire [data_w*6-1:0] v197ibus;
wire [temp_w*6-1:0] v197obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU197 (.l(l[197*data_w +:data_w]), .r(v197ibus), .q(v197obus), .dec(dec[197]));
wire [data_w*6-1:0] v198ibus;
wire [temp_w*6-1:0] v198obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU198 (.l(l[198*data_w +:data_w]), .r(v198ibus), .q(v198obus), .dec(dec[198]));
wire [data_w*6-1:0] v199ibus;
wire [temp_w*6-1:0] v199obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU199 (.l(l[199*data_w +:data_w]), .r(v199ibus), .q(v199obus), .dec(dec[199]));
wire [data_w*6-1:0] v200ibus;
wire [temp_w*6-1:0] v200obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU200 (.l(l[200*data_w +:data_w]), .r(v200ibus), .q(v200obus), .dec(dec[200]));
wire [data_w*6-1:0] v201ibus;
wire [temp_w*6-1:0] v201obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU201 (.l(l[201*data_w +:data_w]), .r(v201ibus), .q(v201obus), .dec(dec[201]));
wire [data_w*6-1:0] v202ibus;
wire [temp_w*6-1:0] v202obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU202 (.l(l[202*data_w +:data_w]), .r(v202ibus), .q(v202obus), .dec(dec[202]));
wire [data_w*6-1:0] v203ibus;
wire [temp_w*6-1:0] v203obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU203 (.l(l[203*data_w +:data_w]), .r(v203ibus), .q(v203obus), .dec(dec[203]));
wire [data_w*6-1:0] v204ibus;
wire [temp_w*6-1:0] v204obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU204 (.l(l[204*data_w +:data_w]), .r(v204ibus), .q(v204obus), .dec(dec[204]));
wire [data_w*6-1:0] v205ibus;
wire [temp_w*6-1:0] v205obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU205 (.l(l[205*data_w +:data_w]), .r(v205ibus), .q(v205obus), .dec(dec[205]));
wire [data_w*6-1:0] v206ibus;
wire [temp_w*6-1:0] v206obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU206 (.l(l[206*data_w +:data_w]), .r(v206ibus), .q(v206obus), .dec(dec[206]));
wire [data_w*6-1:0] v207ibus;
wire [temp_w*6-1:0] v207obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU207 (.l(l[207*data_w +:data_w]), .r(v207ibus), .q(v207obus), .dec(dec[207]));
wire [data_w*6-1:0] v208ibus;
wire [temp_w*6-1:0] v208obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU208 (.l(l[208*data_w +:data_w]), .r(v208ibus), .q(v208obus), .dec(dec[208]));
wire [data_w*6-1:0] v209ibus;
wire [temp_w*6-1:0] v209obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU209 (.l(l[209*data_w +:data_w]), .r(v209ibus), .q(v209obus), .dec(dec[209]));
wire [data_w*6-1:0] v210ibus;
wire [temp_w*6-1:0] v210obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU210 (.l(l[210*data_w +:data_w]), .r(v210ibus), .q(v210obus), .dec(dec[210]));
wire [data_w*6-1:0] v211ibus;
wire [temp_w*6-1:0] v211obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU211 (.l(l[211*data_w +:data_w]), .r(v211ibus), .q(v211obus), .dec(dec[211]));
wire [data_w*6-1:0] v212ibus;
wire [temp_w*6-1:0] v212obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU212 (.l(l[212*data_w +:data_w]), .r(v212ibus), .q(v212obus), .dec(dec[212]));
wire [data_w*6-1:0] v213ibus;
wire [temp_w*6-1:0] v213obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU213 (.l(l[213*data_w +:data_w]), .r(v213ibus), .q(v213obus), .dec(dec[213]));
wire [data_w*6-1:0] v214ibus;
wire [temp_w*6-1:0] v214obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU214 (.l(l[214*data_w +:data_w]), .r(v214ibus), .q(v214obus), .dec(dec[214]));
wire [data_w*6-1:0] v215ibus;
wire [temp_w*6-1:0] v215obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU215 (.l(l[215*data_w +:data_w]), .r(v215ibus), .q(v215obus), .dec(dec[215]));
wire [data_w*6-1:0] v216ibus;
wire [temp_w*6-1:0] v216obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU216 (.l(l[216*data_w +:data_w]), .r(v216ibus), .q(v216obus), .dec(dec[216]));
wire [data_w*6-1:0] v217ibus;
wire [temp_w*6-1:0] v217obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU217 (.l(l[217*data_w +:data_w]), .r(v217ibus), .q(v217obus), .dec(dec[217]));
wire [data_w*6-1:0] v218ibus;
wire [temp_w*6-1:0] v218obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU218 (.l(l[218*data_w +:data_w]), .r(v218ibus), .q(v218obus), .dec(dec[218]));
wire [data_w*6-1:0] v219ibus;
wire [temp_w*6-1:0] v219obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU219 (.l(l[219*data_w +:data_w]), .r(v219ibus), .q(v219obus), .dec(dec[219]));
wire [data_w*6-1:0] v220ibus;
wire [temp_w*6-1:0] v220obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU220 (.l(l[220*data_w +:data_w]), .r(v220ibus), .q(v220obus), .dec(dec[220]));
wire [data_w*6-1:0] v221ibus;
wire [temp_w*6-1:0] v221obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU221 (.l(l[221*data_w +:data_w]), .r(v221ibus), .q(v221obus), .dec(dec[221]));
wire [data_w*6-1:0] v222ibus;
wire [temp_w*6-1:0] v222obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU222 (.l(l[222*data_w +:data_w]), .r(v222ibus), .q(v222obus), .dec(dec[222]));
wire [data_w*6-1:0] v223ibus;
wire [temp_w*6-1:0] v223obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU223 (.l(l[223*data_w +:data_w]), .r(v223ibus), .q(v223obus), .dec(dec[223]));
wire [data_w*6-1:0] v224ibus;
wire [temp_w*6-1:0] v224obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU224 (.l(l[224*data_w +:data_w]), .r(v224ibus), .q(v224obus), .dec(dec[224]));
wire [data_w*6-1:0] v225ibus;
wire [temp_w*6-1:0] v225obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU225 (.l(l[225*data_w +:data_w]), .r(v225ibus), .q(v225obus), .dec(dec[225]));
wire [data_w*6-1:0] v226ibus;
wire [temp_w*6-1:0] v226obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU226 (.l(l[226*data_w +:data_w]), .r(v226ibus), .q(v226obus), .dec(dec[226]));
wire [data_w*6-1:0] v227ibus;
wire [temp_w*6-1:0] v227obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU227 (.l(l[227*data_w +:data_w]), .r(v227ibus), .q(v227obus), .dec(dec[227]));
wire [data_w*6-1:0] v228ibus;
wire [temp_w*6-1:0] v228obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU228 (.l(l[228*data_w +:data_w]), .r(v228ibus), .q(v228obus), .dec(dec[228]));
wire [data_w*6-1:0] v229ibus;
wire [temp_w*6-1:0] v229obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU229 (.l(l[229*data_w +:data_w]), .r(v229ibus), .q(v229obus), .dec(dec[229]));
wire [data_w*6-1:0] v230ibus;
wire [temp_w*6-1:0] v230obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU230 (.l(l[230*data_w +:data_w]), .r(v230ibus), .q(v230obus), .dec(dec[230]));
wire [data_w*6-1:0] v231ibus;
wire [temp_w*6-1:0] v231obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU231 (.l(l[231*data_w +:data_w]), .r(v231ibus), .q(v231obus), .dec(dec[231]));
wire [data_w*6-1:0] v232ibus;
wire [temp_w*6-1:0] v232obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU232 (.l(l[232*data_w +:data_w]), .r(v232ibus), .q(v232obus), .dec(dec[232]));
wire [data_w*6-1:0] v233ibus;
wire [temp_w*6-1:0] v233obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU233 (.l(l[233*data_w +:data_w]), .r(v233ibus), .q(v233obus), .dec(dec[233]));
wire [data_w*6-1:0] v234ibus;
wire [temp_w*6-1:0] v234obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU234 (.l(l[234*data_w +:data_w]), .r(v234ibus), .q(v234obus), .dec(dec[234]));
wire [data_w*6-1:0] v235ibus;
wire [temp_w*6-1:0] v235obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU235 (.l(l[235*data_w +:data_w]), .r(v235ibus), .q(v235obus), .dec(dec[235]));
wire [data_w*6-1:0] v236ibus;
wire [temp_w*6-1:0] v236obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU236 (.l(l[236*data_w +:data_w]), .r(v236ibus), .q(v236obus), .dec(dec[236]));
wire [data_w*6-1:0] v237ibus;
wire [temp_w*6-1:0] v237obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU237 (.l(l[237*data_w +:data_w]), .r(v237ibus), .q(v237obus), .dec(dec[237]));
wire [data_w*6-1:0] v238ibus;
wire [temp_w*6-1:0] v238obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU238 (.l(l[238*data_w +:data_w]), .r(v238ibus), .q(v238obus), .dec(dec[238]));
wire [data_w*6-1:0] v239ibus;
wire [temp_w*6-1:0] v239obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU239 (.l(l[239*data_w +:data_w]), .r(v239ibus), .q(v239obus), .dec(dec[239]));
wire [data_w*6-1:0] v240ibus;
wire [temp_w*6-1:0] v240obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU240 (.l(l[240*data_w +:data_w]), .r(v240ibus), .q(v240obus), .dec(dec[240]));
wire [data_w*6-1:0] v241ibus;
wire [temp_w*6-1:0] v241obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU241 (.l(l[241*data_w +:data_w]), .r(v241ibus), .q(v241obus), .dec(dec[241]));
wire [data_w*6-1:0] v242ibus;
wire [temp_w*6-1:0] v242obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU242 (.l(l[242*data_w +:data_w]), .r(v242ibus), .q(v242obus), .dec(dec[242]));
wire [data_w*6-1:0] v243ibus;
wire [temp_w*6-1:0] v243obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU243 (.l(l[243*data_w +:data_w]), .r(v243ibus), .q(v243obus), .dec(dec[243]));
wire [data_w*6-1:0] v244ibus;
wire [temp_w*6-1:0] v244obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU244 (.l(l[244*data_w +:data_w]), .r(v244ibus), .q(v244obus), .dec(dec[244]));
wire [data_w*6-1:0] v245ibus;
wire [temp_w*6-1:0] v245obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU245 (.l(l[245*data_w +:data_w]), .r(v245ibus), .q(v245obus), .dec(dec[245]));
wire [data_w*6-1:0] v246ibus;
wire [temp_w*6-1:0] v246obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU246 (.l(l[246*data_w +:data_w]), .r(v246ibus), .q(v246obus), .dec(dec[246]));
wire [data_w*6-1:0] v247ibus;
wire [temp_w*6-1:0] v247obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU247 (.l(l[247*data_w +:data_w]), .r(v247ibus), .q(v247obus), .dec(dec[247]));
wire [data_w*6-1:0] v248ibus;
wire [temp_w*6-1:0] v248obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU248 (.l(l[248*data_w +:data_w]), .r(v248ibus), .q(v248obus), .dec(dec[248]));
wire [data_w*6-1:0] v249ibus;
wire [temp_w*6-1:0] v249obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU249 (.l(l[249*data_w +:data_w]), .r(v249ibus), .q(v249obus), .dec(dec[249]));
wire [data_w*6-1:0] v250ibus;
wire [temp_w*6-1:0] v250obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU250 (.l(l[250*data_w +:data_w]), .r(v250ibus), .q(v250obus), .dec(dec[250]));
wire [data_w*6-1:0] v251ibus;
wire [temp_w*6-1:0] v251obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU251 (.l(l[251*data_w +:data_w]), .r(v251ibus), .q(v251obus), .dec(dec[251]));
wire [data_w*6-1:0] v252ibus;
wire [temp_w*6-1:0] v252obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU252 (.l(l[252*data_w +:data_w]), .r(v252ibus), .q(v252obus), .dec(dec[252]));
wire [data_w*6-1:0] v253ibus;
wire [temp_w*6-1:0] v253obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU253 (.l(l[253*data_w +:data_w]), .r(v253ibus), .q(v253obus), .dec(dec[253]));
wire [data_w*6-1:0] v254ibus;
wire [temp_w*6-1:0] v254obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU254 (.l(l[254*data_w +:data_w]), .r(v254ibus), .q(v254obus), .dec(dec[254]));
wire [data_w*6-1:0] v255ibus;
wire [temp_w*6-1:0] v255obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU255 (.l(l[255*data_w +:data_w]), .r(v255ibus), .q(v255obus), .dec(dec[255]));
wire [data_w*6-1:0] v256ibus;
wire [temp_w*6-1:0] v256obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU256 (.l(l[256*data_w +:data_w]), .r(v256ibus), .q(v256obus), .dec(dec[256]));
wire [data_w*6-1:0] v257ibus;
wire [temp_w*6-1:0] v257obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU257 (.l(l[257*data_w +:data_w]), .r(v257ibus), .q(v257obus), .dec(dec[257]));
wire [data_w*6-1:0] v258ibus;
wire [temp_w*6-1:0] v258obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU258 (.l(l[258*data_w +:data_w]), .r(v258ibus), .q(v258obus), .dec(dec[258]));
wire [data_w*6-1:0] v259ibus;
wire [temp_w*6-1:0] v259obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU259 (.l(l[259*data_w +:data_w]), .r(v259ibus), .q(v259obus), .dec(dec[259]));
wire [data_w*6-1:0] v260ibus;
wire [temp_w*6-1:0] v260obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU260 (.l(l[260*data_w +:data_w]), .r(v260ibus), .q(v260obus), .dec(dec[260]));
wire [data_w*6-1:0] v261ibus;
wire [temp_w*6-1:0] v261obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU261 (.l(l[261*data_w +:data_w]), .r(v261ibus), .q(v261obus), .dec(dec[261]));
wire [data_w*6-1:0] v262ibus;
wire [temp_w*6-1:0] v262obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU262 (.l(l[262*data_w +:data_w]), .r(v262ibus), .q(v262obus), .dec(dec[262]));
wire [data_w*6-1:0] v263ibus;
wire [temp_w*6-1:0] v263obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU263 (.l(l[263*data_w +:data_w]), .r(v263ibus), .q(v263obus), .dec(dec[263]));
wire [data_w*6-1:0] v264ibus;
wire [temp_w*6-1:0] v264obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU264 (.l(l[264*data_w +:data_w]), .r(v264ibus), .q(v264obus), .dec(dec[264]));
wire [data_w*6-1:0] v265ibus;
wire [temp_w*6-1:0] v265obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU265 (.l(l[265*data_w +:data_w]), .r(v265ibus), .q(v265obus), .dec(dec[265]));
wire [data_w*6-1:0] v266ibus;
wire [temp_w*6-1:0] v266obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU266 (.l(l[266*data_w +:data_w]), .r(v266ibus), .q(v266obus), .dec(dec[266]));
wire [data_w*6-1:0] v267ibus;
wire [temp_w*6-1:0] v267obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU267 (.l(l[267*data_w +:data_w]), .r(v267ibus), .q(v267obus), .dec(dec[267]));
wire [data_w*6-1:0] v268ibus;
wire [temp_w*6-1:0] v268obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU268 (.l(l[268*data_w +:data_w]), .r(v268ibus), .q(v268obus), .dec(dec[268]));
wire [data_w*6-1:0] v269ibus;
wire [temp_w*6-1:0] v269obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU269 (.l(l[269*data_w +:data_w]), .r(v269ibus), .q(v269obus), .dec(dec[269]));
wire [data_w*6-1:0] v270ibus;
wire [temp_w*6-1:0] v270obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU270 (.l(l[270*data_w +:data_w]), .r(v270ibus), .q(v270obus), .dec(dec[270]));
wire [data_w*6-1:0] v271ibus;
wire [temp_w*6-1:0] v271obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU271 (.l(l[271*data_w +:data_w]), .r(v271ibus), .q(v271obus), .dec(dec[271]));
wire [data_w*6-1:0] v272ibus;
wire [temp_w*6-1:0] v272obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU272 (.l(l[272*data_w +:data_w]), .r(v272ibus), .q(v272obus), .dec(dec[272]));
wire [data_w*6-1:0] v273ibus;
wire [temp_w*6-1:0] v273obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU273 (.l(l[273*data_w +:data_w]), .r(v273ibus), .q(v273obus), .dec(dec[273]));
wire [data_w*6-1:0] v274ibus;
wire [temp_w*6-1:0] v274obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU274 (.l(l[274*data_w +:data_w]), .r(v274ibus), .q(v274obus), .dec(dec[274]));
wire [data_w*6-1:0] v275ibus;
wire [temp_w*6-1:0] v275obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU275 (.l(l[275*data_w +:data_w]), .r(v275ibus), .q(v275obus), .dec(dec[275]));
wire [data_w*6-1:0] v276ibus;
wire [temp_w*6-1:0] v276obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU276 (.l(l[276*data_w +:data_w]), .r(v276ibus), .q(v276obus), .dec(dec[276]));
wire [data_w*6-1:0] v277ibus;
wire [temp_w*6-1:0] v277obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU277 (.l(l[277*data_w +:data_w]), .r(v277ibus), .q(v277obus), .dec(dec[277]));
wire [data_w*6-1:0] v278ibus;
wire [temp_w*6-1:0] v278obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU278 (.l(l[278*data_w +:data_w]), .r(v278ibus), .q(v278obus), .dec(dec[278]));
wire [data_w*6-1:0] v279ibus;
wire [temp_w*6-1:0] v279obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU279 (.l(l[279*data_w +:data_w]), .r(v279ibus), .q(v279obus), .dec(dec[279]));
wire [data_w*6-1:0] v280ibus;
wire [temp_w*6-1:0] v280obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU280 (.l(l[280*data_w +:data_w]), .r(v280ibus), .q(v280obus), .dec(dec[280]));
wire [data_w*6-1:0] v281ibus;
wire [temp_w*6-1:0] v281obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU281 (.l(l[281*data_w +:data_w]), .r(v281ibus), .q(v281obus), .dec(dec[281]));
wire [data_w*6-1:0] v282ibus;
wire [temp_w*6-1:0] v282obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU282 (.l(l[282*data_w +:data_w]), .r(v282ibus), .q(v282obus), .dec(dec[282]));
wire [data_w*6-1:0] v283ibus;
wire [temp_w*6-1:0] v283obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU283 (.l(l[283*data_w +:data_w]), .r(v283ibus), .q(v283obus), .dec(dec[283]));
wire [data_w*6-1:0] v284ibus;
wire [temp_w*6-1:0] v284obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU284 (.l(l[284*data_w +:data_w]), .r(v284ibus), .q(v284obus), .dec(dec[284]));
wire [data_w*6-1:0] v285ibus;
wire [temp_w*6-1:0] v285obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU285 (.l(l[285*data_w +:data_w]), .r(v285ibus), .q(v285obus), .dec(dec[285]));
wire [data_w*6-1:0] v286ibus;
wire [temp_w*6-1:0] v286obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU286 (.l(l[286*data_w +:data_w]), .r(v286ibus), .q(v286obus), .dec(dec[286]));
wire [data_w*6-1:0] v287ibus;
wire [temp_w*6-1:0] v287obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU287 (.l(l[287*data_w +:data_w]), .r(v287ibus), .q(v287obus), .dec(dec[287]));
wire [data_w*3-1:0] v288ibus;
wire [temp_w*3-1:0] v288obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU288 (.l(l[288*data_w +:data_w]), .r(v288ibus), .q(v288obus), .dec(dec[288]));
wire [data_w*3-1:0] v289ibus;
wire [temp_w*3-1:0] v289obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU289 (.l(l[289*data_w +:data_w]), .r(v289ibus), .q(v289obus), .dec(dec[289]));
wire [data_w*3-1:0] v290ibus;
wire [temp_w*3-1:0] v290obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU290 (.l(l[290*data_w +:data_w]), .r(v290ibus), .q(v290obus), .dec(dec[290]));
wire [data_w*3-1:0] v291ibus;
wire [temp_w*3-1:0] v291obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU291 (.l(l[291*data_w +:data_w]), .r(v291ibus), .q(v291obus), .dec(dec[291]));
wire [data_w*3-1:0] v292ibus;
wire [temp_w*3-1:0] v292obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU292 (.l(l[292*data_w +:data_w]), .r(v292ibus), .q(v292obus), .dec(dec[292]));
wire [data_w*3-1:0] v293ibus;
wire [temp_w*3-1:0] v293obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU293 (.l(l[293*data_w +:data_w]), .r(v293ibus), .q(v293obus), .dec(dec[293]));
wire [data_w*3-1:0] v294ibus;
wire [temp_w*3-1:0] v294obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU294 (.l(l[294*data_w +:data_w]), .r(v294ibus), .q(v294obus), .dec(dec[294]));
wire [data_w*3-1:0] v295ibus;
wire [temp_w*3-1:0] v295obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU295 (.l(l[295*data_w +:data_w]), .r(v295ibus), .q(v295obus), .dec(dec[295]));
wire [data_w*3-1:0] v296ibus;
wire [temp_w*3-1:0] v296obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU296 (.l(l[296*data_w +:data_w]), .r(v296ibus), .q(v296obus), .dec(dec[296]));
wire [data_w*3-1:0] v297ibus;
wire [temp_w*3-1:0] v297obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU297 (.l(l[297*data_w +:data_w]), .r(v297ibus), .q(v297obus), .dec(dec[297]));
wire [data_w*3-1:0] v298ibus;
wire [temp_w*3-1:0] v298obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU298 (.l(l[298*data_w +:data_w]), .r(v298ibus), .q(v298obus), .dec(dec[298]));
wire [data_w*3-1:0] v299ibus;
wire [temp_w*3-1:0] v299obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU299 (.l(l[299*data_w +:data_w]), .r(v299ibus), .q(v299obus), .dec(dec[299]));
wire [data_w*3-1:0] v300ibus;
wire [temp_w*3-1:0] v300obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU300 (.l(l[300*data_w +:data_w]), .r(v300ibus), .q(v300obus), .dec(dec[300]));
wire [data_w*3-1:0] v301ibus;
wire [temp_w*3-1:0] v301obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU301 (.l(l[301*data_w +:data_w]), .r(v301ibus), .q(v301obus), .dec(dec[301]));
wire [data_w*3-1:0] v302ibus;
wire [temp_w*3-1:0] v302obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU302 (.l(l[302*data_w +:data_w]), .r(v302ibus), .q(v302obus), .dec(dec[302]));
wire [data_w*3-1:0] v303ibus;
wire [temp_w*3-1:0] v303obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU303 (.l(l[303*data_w +:data_w]), .r(v303ibus), .q(v303obus), .dec(dec[303]));
wire [data_w*3-1:0] v304ibus;
wire [temp_w*3-1:0] v304obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU304 (.l(l[304*data_w +:data_w]), .r(v304ibus), .q(v304obus), .dec(dec[304]));
wire [data_w*3-1:0] v305ibus;
wire [temp_w*3-1:0] v305obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU305 (.l(l[305*data_w +:data_w]), .r(v305ibus), .q(v305obus), .dec(dec[305]));
wire [data_w*3-1:0] v306ibus;
wire [temp_w*3-1:0] v306obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU306 (.l(l[306*data_w +:data_w]), .r(v306ibus), .q(v306obus), .dec(dec[306]));
wire [data_w*3-1:0] v307ibus;
wire [temp_w*3-1:0] v307obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU307 (.l(l[307*data_w +:data_w]), .r(v307ibus), .q(v307obus), .dec(dec[307]));
wire [data_w*3-1:0] v308ibus;
wire [temp_w*3-1:0] v308obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU308 (.l(l[308*data_w +:data_w]), .r(v308ibus), .q(v308obus), .dec(dec[308]));
wire [data_w*3-1:0] v309ibus;
wire [temp_w*3-1:0] v309obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU309 (.l(l[309*data_w +:data_w]), .r(v309ibus), .q(v309obus), .dec(dec[309]));
wire [data_w*3-1:0] v310ibus;
wire [temp_w*3-1:0] v310obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU310 (.l(l[310*data_w +:data_w]), .r(v310ibus), .q(v310obus), .dec(dec[310]));
wire [data_w*3-1:0] v311ibus;
wire [temp_w*3-1:0] v311obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU311 (.l(l[311*data_w +:data_w]), .r(v311ibus), .q(v311obus), .dec(dec[311]));
wire [data_w*3-1:0] v312ibus;
wire [temp_w*3-1:0] v312obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU312 (.l(l[312*data_w +:data_w]), .r(v312ibus), .q(v312obus), .dec(dec[312]));
wire [data_w*3-1:0] v313ibus;
wire [temp_w*3-1:0] v313obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU313 (.l(l[313*data_w +:data_w]), .r(v313ibus), .q(v313obus), .dec(dec[313]));
wire [data_w*3-1:0] v314ibus;
wire [temp_w*3-1:0] v314obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU314 (.l(l[314*data_w +:data_w]), .r(v314ibus), .q(v314obus), .dec(dec[314]));
wire [data_w*3-1:0] v315ibus;
wire [temp_w*3-1:0] v315obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU315 (.l(l[315*data_w +:data_w]), .r(v315ibus), .q(v315obus), .dec(dec[315]));
wire [data_w*3-1:0] v316ibus;
wire [temp_w*3-1:0] v316obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU316 (.l(l[316*data_w +:data_w]), .r(v316ibus), .q(v316obus), .dec(dec[316]));
wire [data_w*3-1:0] v317ibus;
wire [temp_w*3-1:0] v317obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU317 (.l(l[317*data_w +:data_w]), .r(v317ibus), .q(v317obus), .dec(dec[317]));
wire [data_w*3-1:0] v318ibus;
wire [temp_w*3-1:0] v318obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU318 (.l(l[318*data_w +:data_w]), .r(v318ibus), .q(v318obus), .dec(dec[318]));
wire [data_w*3-1:0] v319ibus;
wire [temp_w*3-1:0] v319obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU319 (.l(l[319*data_w +:data_w]), .r(v319ibus), .q(v319obus), .dec(dec[319]));
wire [data_w*3-1:0] v320ibus;
wire [temp_w*3-1:0] v320obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU320 (.l(l[320*data_w +:data_w]), .r(v320ibus), .q(v320obus), .dec(dec[320]));
wire [data_w*3-1:0] v321ibus;
wire [temp_w*3-1:0] v321obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU321 (.l(l[321*data_w +:data_w]), .r(v321ibus), .q(v321obus), .dec(dec[321]));
wire [data_w*3-1:0] v322ibus;
wire [temp_w*3-1:0] v322obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU322 (.l(l[322*data_w +:data_w]), .r(v322ibus), .q(v322obus), .dec(dec[322]));
wire [data_w*3-1:0] v323ibus;
wire [temp_w*3-1:0] v323obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU323 (.l(l[323*data_w +:data_w]), .r(v323ibus), .q(v323obus), .dec(dec[323]));
wire [data_w*3-1:0] v324ibus;
wire [temp_w*3-1:0] v324obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU324 (.l(l[324*data_w +:data_w]), .r(v324ibus), .q(v324obus), .dec(dec[324]));
wire [data_w*3-1:0] v325ibus;
wire [temp_w*3-1:0] v325obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU325 (.l(l[325*data_w +:data_w]), .r(v325ibus), .q(v325obus), .dec(dec[325]));
wire [data_w*3-1:0] v326ibus;
wire [temp_w*3-1:0] v326obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU326 (.l(l[326*data_w +:data_w]), .r(v326ibus), .q(v326obus), .dec(dec[326]));
wire [data_w*3-1:0] v327ibus;
wire [temp_w*3-1:0] v327obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU327 (.l(l[327*data_w +:data_w]), .r(v327ibus), .q(v327obus), .dec(dec[327]));
wire [data_w*3-1:0] v328ibus;
wire [temp_w*3-1:0] v328obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU328 (.l(l[328*data_w +:data_w]), .r(v328ibus), .q(v328obus), .dec(dec[328]));
wire [data_w*3-1:0] v329ibus;
wire [temp_w*3-1:0] v329obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU329 (.l(l[329*data_w +:data_w]), .r(v329ibus), .q(v329obus), .dec(dec[329]));
wire [data_w*3-1:0] v330ibus;
wire [temp_w*3-1:0] v330obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU330 (.l(l[330*data_w +:data_w]), .r(v330ibus), .q(v330obus), .dec(dec[330]));
wire [data_w*3-1:0] v331ibus;
wire [temp_w*3-1:0] v331obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU331 (.l(l[331*data_w +:data_w]), .r(v331ibus), .q(v331obus), .dec(dec[331]));
wire [data_w*3-1:0] v332ibus;
wire [temp_w*3-1:0] v332obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU332 (.l(l[332*data_w +:data_w]), .r(v332ibus), .q(v332obus), .dec(dec[332]));
wire [data_w*3-1:0] v333ibus;
wire [temp_w*3-1:0] v333obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU333 (.l(l[333*data_w +:data_w]), .r(v333ibus), .q(v333obus), .dec(dec[333]));
wire [data_w*3-1:0] v334ibus;
wire [temp_w*3-1:0] v334obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU334 (.l(l[334*data_w +:data_w]), .r(v334ibus), .q(v334obus), .dec(dec[334]));
wire [data_w*3-1:0] v335ibus;
wire [temp_w*3-1:0] v335obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU335 (.l(l[335*data_w +:data_w]), .r(v335ibus), .q(v335obus), .dec(dec[335]));
wire [data_w*3-1:0] v336ibus;
wire [temp_w*3-1:0] v336obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU336 (.l(l[336*data_w +:data_w]), .r(v336ibus), .q(v336obus), .dec(dec[336]));
wire [data_w*3-1:0] v337ibus;
wire [temp_w*3-1:0] v337obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU337 (.l(l[337*data_w +:data_w]), .r(v337ibus), .q(v337obus), .dec(dec[337]));
wire [data_w*3-1:0] v338ibus;
wire [temp_w*3-1:0] v338obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU338 (.l(l[338*data_w +:data_w]), .r(v338ibus), .q(v338obus), .dec(dec[338]));
wire [data_w*3-1:0] v339ibus;
wire [temp_w*3-1:0] v339obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU339 (.l(l[339*data_w +:data_w]), .r(v339ibus), .q(v339obus), .dec(dec[339]));
wire [data_w*3-1:0] v340ibus;
wire [temp_w*3-1:0] v340obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU340 (.l(l[340*data_w +:data_w]), .r(v340ibus), .q(v340obus), .dec(dec[340]));
wire [data_w*3-1:0] v341ibus;
wire [temp_w*3-1:0] v341obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU341 (.l(l[341*data_w +:data_w]), .r(v341ibus), .q(v341obus), .dec(dec[341]));
wire [data_w*3-1:0] v342ibus;
wire [temp_w*3-1:0] v342obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU342 (.l(l[342*data_w +:data_w]), .r(v342ibus), .q(v342obus), .dec(dec[342]));
wire [data_w*3-1:0] v343ibus;
wire [temp_w*3-1:0] v343obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU343 (.l(l[343*data_w +:data_w]), .r(v343ibus), .q(v343obus), .dec(dec[343]));
wire [data_w*3-1:0] v344ibus;
wire [temp_w*3-1:0] v344obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU344 (.l(l[344*data_w +:data_w]), .r(v344ibus), .q(v344obus), .dec(dec[344]));
wire [data_w*3-1:0] v345ibus;
wire [temp_w*3-1:0] v345obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU345 (.l(l[345*data_w +:data_w]), .r(v345ibus), .q(v345obus), .dec(dec[345]));
wire [data_w*3-1:0] v346ibus;
wire [temp_w*3-1:0] v346obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU346 (.l(l[346*data_w +:data_w]), .r(v346ibus), .q(v346obus), .dec(dec[346]));
wire [data_w*3-1:0] v347ibus;
wire [temp_w*3-1:0] v347obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU347 (.l(l[347*data_w +:data_w]), .r(v347ibus), .q(v347obus), .dec(dec[347]));
wire [data_w*3-1:0] v348ibus;
wire [temp_w*3-1:0] v348obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU348 (.l(l[348*data_w +:data_w]), .r(v348ibus), .q(v348obus), .dec(dec[348]));
wire [data_w*3-1:0] v349ibus;
wire [temp_w*3-1:0] v349obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU349 (.l(l[349*data_w +:data_w]), .r(v349ibus), .q(v349obus), .dec(dec[349]));
wire [data_w*3-1:0] v350ibus;
wire [temp_w*3-1:0] v350obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU350 (.l(l[350*data_w +:data_w]), .r(v350ibus), .q(v350obus), .dec(dec[350]));
wire [data_w*3-1:0] v351ibus;
wire [temp_w*3-1:0] v351obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU351 (.l(l[351*data_w +:data_w]), .r(v351ibus), .q(v351obus), .dec(dec[351]));
wire [data_w*3-1:0] v352ibus;
wire [temp_w*3-1:0] v352obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU352 (.l(l[352*data_w +:data_w]), .r(v352ibus), .q(v352obus), .dec(dec[352]));
wire [data_w*3-1:0] v353ibus;
wire [temp_w*3-1:0] v353obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU353 (.l(l[353*data_w +:data_w]), .r(v353ibus), .q(v353obus), .dec(dec[353]));
wire [data_w*3-1:0] v354ibus;
wire [temp_w*3-1:0] v354obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU354 (.l(l[354*data_w +:data_w]), .r(v354ibus), .q(v354obus), .dec(dec[354]));
wire [data_w*3-1:0] v355ibus;
wire [temp_w*3-1:0] v355obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU355 (.l(l[355*data_w +:data_w]), .r(v355ibus), .q(v355obus), .dec(dec[355]));
wire [data_w*3-1:0] v356ibus;
wire [temp_w*3-1:0] v356obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU356 (.l(l[356*data_w +:data_w]), .r(v356ibus), .q(v356obus), .dec(dec[356]));
wire [data_w*3-1:0] v357ibus;
wire [temp_w*3-1:0] v357obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU357 (.l(l[357*data_w +:data_w]), .r(v357ibus), .q(v357obus), .dec(dec[357]));
wire [data_w*3-1:0] v358ibus;
wire [temp_w*3-1:0] v358obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU358 (.l(l[358*data_w +:data_w]), .r(v358ibus), .q(v358obus), .dec(dec[358]));
wire [data_w*3-1:0] v359ibus;
wire [temp_w*3-1:0] v359obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU359 (.l(l[359*data_w +:data_w]), .r(v359ibus), .q(v359obus), .dec(dec[359]));
wire [data_w*3-1:0] v360ibus;
wire [temp_w*3-1:0] v360obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU360 (.l(l[360*data_w +:data_w]), .r(v360ibus), .q(v360obus), .dec(dec[360]));
wire [data_w*3-1:0] v361ibus;
wire [temp_w*3-1:0] v361obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU361 (.l(l[361*data_w +:data_w]), .r(v361ibus), .q(v361obus), .dec(dec[361]));
wire [data_w*3-1:0] v362ibus;
wire [temp_w*3-1:0] v362obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU362 (.l(l[362*data_w +:data_w]), .r(v362ibus), .q(v362obus), .dec(dec[362]));
wire [data_w*3-1:0] v363ibus;
wire [temp_w*3-1:0] v363obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU363 (.l(l[363*data_w +:data_w]), .r(v363ibus), .q(v363obus), .dec(dec[363]));
wire [data_w*3-1:0] v364ibus;
wire [temp_w*3-1:0] v364obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU364 (.l(l[364*data_w +:data_w]), .r(v364ibus), .q(v364obus), .dec(dec[364]));
wire [data_w*3-1:0] v365ibus;
wire [temp_w*3-1:0] v365obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU365 (.l(l[365*data_w +:data_w]), .r(v365ibus), .q(v365obus), .dec(dec[365]));
wire [data_w*3-1:0] v366ibus;
wire [temp_w*3-1:0] v366obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU366 (.l(l[366*data_w +:data_w]), .r(v366ibus), .q(v366obus), .dec(dec[366]));
wire [data_w*3-1:0] v367ibus;
wire [temp_w*3-1:0] v367obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU367 (.l(l[367*data_w +:data_w]), .r(v367ibus), .q(v367obus), .dec(dec[367]));
wire [data_w*3-1:0] v368ibus;
wire [temp_w*3-1:0] v368obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU368 (.l(l[368*data_w +:data_w]), .r(v368ibus), .q(v368obus), .dec(dec[368]));
wire [data_w*3-1:0] v369ibus;
wire [temp_w*3-1:0] v369obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU369 (.l(l[369*data_w +:data_w]), .r(v369ibus), .q(v369obus), .dec(dec[369]));
wire [data_w*3-1:0] v370ibus;
wire [temp_w*3-1:0] v370obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU370 (.l(l[370*data_w +:data_w]), .r(v370ibus), .q(v370obus), .dec(dec[370]));
wire [data_w*3-1:0] v371ibus;
wire [temp_w*3-1:0] v371obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU371 (.l(l[371*data_w +:data_w]), .r(v371ibus), .q(v371obus), .dec(dec[371]));
wire [data_w*3-1:0] v372ibus;
wire [temp_w*3-1:0] v372obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU372 (.l(l[372*data_w +:data_w]), .r(v372ibus), .q(v372obus), .dec(dec[372]));
wire [data_w*3-1:0] v373ibus;
wire [temp_w*3-1:0] v373obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU373 (.l(l[373*data_w +:data_w]), .r(v373ibus), .q(v373obus), .dec(dec[373]));
wire [data_w*3-1:0] v374ibus;
wire [temp_w*3-1:0] v374obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU374 (.l(l[374*data_w +:data_w]), .r(v374ibus), .q(v374obus), .dec(dec[374]));
wire [data_w*3-1:0] v375ibus;
wire [temp_w*3-1:0] v375obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU375 (.l(l[375*data_w +:data_w]), .r(v375ibus), .q(v375obus), .dec(dec[375]));
wire [data_w*3-1:0] v376ibus;
wire [temp_w*3-1:0] v376obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU376 (.l(l[376*data_w +:data_w]), .r(v376ibus), .q(v376obus), .dec(dec[376]));
wire [data_w*3-1:0] v377ibus;
wire [temp_w*3-1:0] v377obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU377 (.l(l[377*data_w +:data_w]), .r(v377ibus), .q(v377obus), .dec(dec[377]));
wire [data_w*3-1:0] v378ibus;
wire [temp_w*3-1:0] v378obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU378 (.l(l[378*data_w +:data_w]), .r(v378ibus), .q(v378obus), .dec(dec[378]));
wire [data_w*3-1:0] v379ibus;
wire [temp_w*3-1:0] v379obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU379 (.l(l[379*data_w +:data_w]), .r(v379ibus), .q(v379obus), .dec(dec[379]));
wire [data_w*3-1:0] v380ibus;
wire [temp_w*3-1:0] v380obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU380 (.l(l[380*data_w +:data_w]), .r(v380ibus), .q(v380obus), .dec(dec[380]));
wire [data_w*3-1:0] v381ibus;
wire [temp_w*3-1:0] v381obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU381 (.l(l[381*data_w +:data_w]), .r(v381ibus), .q(v381obus), .dec(dec[381]));
wire [data_w*3-1:0] v382ibus;
wire [temp_w*3-1:0] v382obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU382 (.l(l[382*data_w +:data_w]), .r(v382ibus), .q(v382obus), .dec(dec[382]));
wire [data_w*3-1:0] v383ibus;
wire [temp_w*3-1:0] v383obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU383 (.l(l[383*data_w +:data_w]), .r(v383ibus), .q(v383obus), .dec(dec[383]));
wire [data_w*3-1:0] v384ibus;
wire [temp_w*3-1:0] v384obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU384 (.l(l[384*data_w +:data_w]), .r(v384ibus), .q(v384obus), .dec(dec[384]));
wire [data_w*3-1:0] v385ibus;
wire [temp_w*3-1:0] v385obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU385 (.l(l[385*data_w +:data_w]), .r(v385ibus), .q(v385obus), .dec(dec[385]));
wire [data_w*3-1:0] v386ibus;
wire [temp_w*3-1:0] v386obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU386 (.l(l[386*data_w +:data_w]), .r(v386ibus), .q(v386obus), .dec(dec[386]));
wire [data_w*3-1:0] v387ibus;
wire [temp_w*3-1:0] v387obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU387 (.l(l[387*data_w +:data_w]), .r(v387ibus), .q(v387obus), .dec(dec[387]));
wire [data_w*3-1:0] v388ibus;
wire [temp_w*3-1:0] v388obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU388 (.l(l[388*data_w +:data_w]), .r(v388ibus), .q(v388obus), .dec(dec[388]));
wire [data_w*3-1:0] v389ibus;
wire [temp_w*3-1:0] v389obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU389 (.l(l[389*data_w +:data_w]), .r(v389ibus), .q(v389obus), .dec(dec[389]));
wire [data_w*3-1:0] v390ibus;
wire [temp_w*3-1:0] v390obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU390 (.l(l[390*data_w +:data_w]), .r(v390ibus), .q(v390obus), .dec(dec[390]));
wire [data_w*3-1:0] v391ibus;
wire [temp_w*3-1:0] v391obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU391 (.l(l[391*data_w +:data_w]), .r(v391ibus), .q(v391obus), .dec(dec[391]));
wire [data_w*3-1:0] v392ibus;
wire [temp_w*3-1:0] v392obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU392 (.l(l[392*data_w +:data_w]), .r(v392ibus), .q(v392obus), .dec(dec[392]));
wire [data_w*3-1:0] v393ibus;
wire [temp_w*3-1:0] v393obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU393 (.l(l[393*data_w +:data_w]), .r(v393ibus), .q(v393obus), .dec(dec[393]));
wire [data_w*3-1:0] v394ibus;
wire [temp_w*3-1:0] v394obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU394 (.l(l[394*data_w +:data_w]), .r(v394ibus), .q(v394obus), .dec(dec[394]));
wire [data_w*3-1:0] v395ibus;
wire [temp_w*3-1:0] v395obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU395 (.l(l[395*data_w +:data_w]), .r(v395ibus), .q(v395obus), .dec(dec[395]));
wire [data_w*3-1:0] v396ibus;
wire [temp_w*3-1:0] v396obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU396 (.l(l[396*data_w +:data_w]), .r(v396ibus), .q(v396obus), .dec(dec[396]));
wire [data_w*3-1:0] v397ibus;
wire [temp_w*3-1:0] v397obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU397 (.l(l[397*data_w +:data_w]), .r(v397ibus), .q(v397obus), .dec(dec[397]));
wire [data_w*3-1:0] v398ibus;
wire [temp_w*3-1:0] v398obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU398 (.l(l[398*data_w +:data_w]), .r(v398ibus), .q(v398obus), .dec(dec[398]));
wire [data_w*3-1:0] v399ibus;
wire [temp_w*3-1:0] v399obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU399 (.l(l[399*data_w +:data_w]), .r(v399ibus), .q(v399obus), .dec(dec[399]));
wire [data_w*3-1:0] v400ibus;
wire [temp_w*3-1:0] v400obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU400 (.l(l[400*data_w +:data_w]), .r(v400ibus), .q(v400obus), .dec(dec[400]));
wire [data_w*3-1:0] v401ibus;
wire [temp_w*3-1:0] v401obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU401 (.l(l[401*data_w +:data_w]), .r(v401ibus), .q(v401obus), .dec(dec[401]));
wire [data_w*3-1:0] v402ibus;
wire [temp_w*3-1:0] v402obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU402 (.l(l[402*data_w +:data_w]), .r(v402ibus), .q(v402obus), .dec(dec[402]));
wire [data_w*3-1:0] v403ibus;
wire [temp_w*3-1:0] v403obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU403 (.l(l[403*data_w +:data_w]), .r(v403ibus), .q(v403obus), .dec(dec[403]));
wire [data_w*3-1:0] v404ibus;
wire [temp_w*3-1:0] v404obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU404 (.l(l[404*data_w +:data_w]), .r(v404ibus), .q(v404obus), .dec(dec[404]));
wire [data_w*3-1:0] v405ibus;
wire [temp_w*3-1:0] v405obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU405 (.l(l[405*data_w +:data_w]), .r(v405ibus), .q(v405obus), .dec(dec[405]));
wire [data_w*3-1:0] v406ibus;
wire [temp_w*3-1:0] v406obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU406 (.l(l[406*data_w +:data_w]), .r(v406ibus), .q(v406obus), .dec(dec[406]));
wire [data_w*3-1:0] v407ibus;
wire [temp_w*3-1:0] v407obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU407 (.l(l[407*data_w +:data_w]), .r(v407ibus), .q(v407obus), .dec(dec[407]));
wire [data_w*3-1:0] v408ibus;
wire [temp_w*3-1:0] v408obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU408 (.l(l[408*data_w +:data_w]), .r(v408ibus), .q(v408obus), .dec(dec[408]));
wire [data_w*3-1:0] v409ibus;
wire [temp_w*3-1:0] v409obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU409 (.l(l[409*data_w +:data_w]), .r(v409ibus), .q(v409obus), .dec(dec[409]));
wire [data_w*3-1:0] v410ibus;
wire [temp_w*3-1:0] v410obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU410 (.l(l[410*data_w +:data_w]), .r(v410ibus), .q(v410obus), .dec(dec[410]));
wire [data_w*3-1:0] v411ibus;
wire [temp_w*3-1:0] v411obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU411 (.l(l[411*data_w +:data_w]), .r(v411ibus), .q(v411obus), .dec(dec[411]));
wire [data_w*3-1:0] v412ibus;
wire [temp_w*3-1:0] v412obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU412 (.l(l[412*data_w +:data_w]), .r(v412ibus), .q(v412obus), .dec(dec[412]));
wire [data_w*3-1:0] v413ibus;
wire [temp_w*3-1:0] v413obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU413 (.l(l[413*data_w +:data_w]), .r(v413ibus), .q(v413obus), .dec(dec[413]));
wire [data_w*3-1:0] v414ibus;
wire [temp_w*3-1:0] v414obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU414 (.l(l[414*data_w +:data_w]), .r(v414ibus), .q(v414obus), .dec(dec[414]));
wire [data_w*3-1:0] v415ibus;
wire [temp_w*3-1:0] v415obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU415 (.l(l[415*data_w +:data_w]), .r(v415ibus), .q(v415obus), .dec(dec[415]));
wire [data_w*3-1:0] v416ibus;
wire [temp_w*3-1:0] v416obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU416 (.l(l[416*data_w +:data_w]), .r(v416ibus), .q(v416obus), .dec(dec[416]));
wire [data_w*3-1:0] v417ibus;
wire [temp_w*3-1:0] v417obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU417 (.l(l[417*data_w +:data_w]), .r(v417ibus), .q(v417obus), .dec(dec[417]));
wire [data_w*3-1:0] v418ibus;
wire [temp_w*3-1:0] v418obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU418 (.l(l[418*data_w +:data_w]), .r(v418ibus), .q(v418obus), .dec(dec[418]));
wire [data_w*3-1:0] v419ibus;
wire [temp_w*3-1:0] v419obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU419 (.l(l[419*data_w +:data_w]), .r(v419ibus), .q(v419obus), .dec(dec[419]));
wire [data_w*3-1:0] v420ibus;
wire [temp_w*3-1:0] v420obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU420 (.l(l[420*data_w +:data_w]), .r(v420ibus), .q(v420obus), .dec(dec[420]));
wire [data_w*3-1:0] v421ibus;
wire [temp_w*3-1:0] v421obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU421 (.l(l[421*data_w +:data_w]), .r(v421ibus), .q(v421obus), .dec(dec[421]));
wire [data_w*3-1:0] v422ibus;
wire [temp_w*3-1:0] v422obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU422 (.l(l[422*data_w +:data_w]), .r(v422ibus), .q(v422obus), .dec(dec[422]));
wire [data_w*3-1:0] v423ibus;
wire [temp_w*3-1:0] v423obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU423 (.l(l[423*data_w +:data_w]), .r(v423ibus), .q(v423obus), .dec(dec[423]));
wire [data_w*3-1:0] v424ibus;
wire [temp_w*3-1:0] v424obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU424 (.l(l[424*data_w +:data_w]), .r(v424ibus), .q(v424obus), .dec(dec[424]));
wire [data_w*3-1:0] v425ibus;
wire [temp_w*3-1:0] v425obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU425 (.l(l[425*data_w +:data_w]), .r(v425ibus), .q(v425obus), .dec(dec[425]));
wire [data_w*3-1:0] v426ibus;
wire [temp_w*3-1:0] v426obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU426 (.l(l[426*data_w +:data_w]), .r(v426ibus), .q(v426obus), .dec(dec[426]));
wire [data_w*3-1:0] v427ibus;
wire [temp_w*3-1:0] v427obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU427 (.l(l[427*data_w +:data_w]), .r(v427ibus), .q(v427obus), .dec(dec[427]));
wire [data_w*3-1:0] v428ibus;
wire [temp_w*3-1:0] v428obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU428 (.l(l[428*data_w +:data_w]), .r(v428ibus), .q(v428obus), .dec(dec[428]));
wire [data_w*3-1:0] v429ibus;
wire [temp_w*3-1:0] v429obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU429 (.l(l[429*data_w +:data_w]), .r(v429ibus), .q(v429obus), .dec(dec[429]));
wire [data_w*3-1:0] v430ibus;
wire [temp_w*3-1:0] v430obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU430 (.l(l[430*data_w +:data_w]), .r(v430ibus), .q(v430obus), .dec(dec[430]));
wire [data_w*3-1:0] v431ibus;
wire [temp_w*3-1:0] v431obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU431 (.l(l[431*data_w +:data_w]), .r(v431ibus), .q(v431obus), .dec(dec[431]));
wire [data_w*3-1:0] v432ibus;
wire [temp_w*3-1:0] v432obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU432 (.l(l[432*data_w +:data_w]), .r(v432ibus), .q(v432obus), .dec(dec[432]));
wire [data_w*3-1:0] v433ibus;
wire [temp_w*3-1:0] v433obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU433 (.l(l[433*data_w +:data_w]), .r(v433ibus), .q(v433obus), .dec(dec[433]));
wire [data_w*3-1:0] v434ibus;
wire [temp_w*3-1:0] v434obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU434 (.l(l[434*data_w +:data_w]), .r(v434ibus), .q(v434obus), .dec(dec[434]));
wire [data_w*3-1:0] v435ibus;
wire [temp_w*3-1:0] v435obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU435 (.l(l[435*data_w +:data_w]), .r(v435ibus), .q(v435obus), .dec(dec[435]));
wire [data_w*3-1:0] v436ibus;
wire [temp_w*3-1:0] v436obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU436 (.l(l[436*data_w +:data_w]), .r(v436ibus), .q(v436obus), .dec(dec[436]));
wire [data_w*3-1:0] v437ibus;
wire [temp_w*3-1:0] v437obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU437 (.l(l[437*data_w +:data_w]), .r(v437ibus), .q(v437obus), .dec(dec[437]));
wire [data_w*3-1:0] v438ibus;
wire [temp_w*3-1:0] v438obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU438 (.l(l[438*data_w +:data_w]), .r(v438ibus), .q(v438obus), .dec(dec[438]));
wire [data_w*3-1:0] v439ibus;
wire [temp_w*3-1:0] v439obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU439 (.l(l[439*data_w +:data_w]), .r(v439ibus), .q(v439obus), .dec(dec[439]));
wire [data_w*3-1:0] v440ibus;
wire [temp_w*3-1:0] v440obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU440 (.l(l[440*data_w +:data_w]), .r(v440ibus), .q(v440obus), .dec(dec[440]));
wire [data_w*3-1:0] v441ibus;
wire [temp_w*3-1:0] v441obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU441 (.l(l[441*data_w +:data_w]), .r(v441ibus), .q(v441obus), .dec(dec[441]));
wire [data_w*3-1:0] v442ibus;
wire [temp_w*3-1:0] v442obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU442 (.l(l[442*data_w +:data_w]), .r(v442ibus), .q(v442obus), .dec(dec[442]));
wire [data_w*3-1:0] v443ibus;
wire [temp_w*3-1:0] v443obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU443 (.l(l[443*data_w +:data_w]), .r(v443ibus), .q(v443obus), .dec(dec[443]));
wire [data_w*3-1:0] v444ibus;
wire [temp_w*3-1:0] v444obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU444 (.l(l[444*data_w +:data_w]), .r(v444ibus), .q(v444obus), .dec(dec[444]));
wire [data_w*3-1:0] v445ibus;
wire [temp_w*3-1:0] v445obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU445 (.l(l[445*data_w +:data_w]), .r(v445ibus), .q(v445obus), .dec(dec[445]));
wire [data_w*3-1:0] v446ibus;
wire [temp_w*3-1:0] v446obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU446 (.l(l[446*data_w +:data_w]), .r(v446ibus), .q(v446obus), .dec(dec[446]));
wire [data_w*3-1:0] v447ibus;
wire [temp_w*3-1:0] v447obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU447 (.l(l[447*data_w +:data_w]), .r(v447ibus), .q(v447obus), .dec(dec[447]));
wire [data_w*3-1:0] v448ibus;
wire [temp_w*3-1:0] v448obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU448 (.l(l[448*data_w +:data_w]), .r(v448ibus), .q(v448obus), .dec(dec[448]));
wire [data_w*3-1:0] v449ibus;
wire [temp_w*3-1:0] v449obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU449 (.l(l[449*data_w +:data_w]), .r(v449ibus), .q(v449obus), .dec(dec[449]));
wire [data_w*3-1:0] v450ibus;
wire [temp_w*3-1:0] v450obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU450 (.l(l[450*data_w +:data_w]), .r(v450ibus), .q(v450obus), .dec(dec[450]));
wire [data_w*3-1:0] v451ibus;
wire [temp_w*3-1:0] v451obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU451 (.l(l[451*data_w +:data_w]), .r(v451ibus), .q(v451obus), .dec(dec[451]));
wire [data_w*3-1:0] v452ibus;
wire [temp_w*3-1:0] v452obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU452 (.l(l[452*data_w +:data_w]), .r(v452ibus), .q(v452obus), .dec(dec[452]));
wire [data_w*3-1:0] v453ibus;
wire [temp_w*3-1:0] v453obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU453 (.l(l[453*data_w +:data_w]), .r(v453ibus), .q(v453obus), .dec(dec[453]));
wire [data_w*3-1:0] v454ibus;
wire [temp_w*3-1:0] v454obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU454 (.l(l[454*data_w +:data_w]), .r(v454ibus), .q(v454obus), .dec(dec[454]));
wire [data_w*3-1:0] v455ibus;
wire [temp_w*3-1:0] v455obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU455 (.l(l[455*data_w +:data_w]), .r(v455ibus), .q(v455obus), .dec(dec[455]));
wire [data_w*3-1:0] v456ibus;
wire [temp_w*3-1:0] v456obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU456 (.l(l[456*data_w +:data_w]), .r(v456ibus), .q(v456obus), .dec(dec[456]));
wire [data_w*3-1:0] v457ibus;
wire [temp_w*3-1:0] v457obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU457 (.l(l[457*data_w +:data_w]), .r(v457ibus), .q(v457obus), .dec(dec[457]));
wire [data_w*3-1:0] v458ibus;
wire [temp_w*3-1:0] v458obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU458 (.l(l[458*data_w +:data_w]), .r(v458ibus), .q(v458obus), .dec(dec[458]));
wire [data_w*3-1:0] v459ibus;
wire [temp_w*3-1:0] v459obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU459 (.l(l[459*data_w +:data_w]), .r(v459ibus), .q(v459obus), .dec(dec[459]));
wire [data_w*3-1:0] v460ibus;
wire [temp_w*3-1:0] v460obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU460 (.l(l[460*data_w +:data_w]), .r(v460ibus), .q(v460obus), .dec(dec[460]));
wire [data_w*3-1:0] v461ibus;
wire [temp_w*3-1:0] v461obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU461 (.l(l[461*data_w +:data_w]), .r(v461ibus), .q(v461obus), .dec(dec[461]));
wire [data_w*3-1:0] v462ibus;
wire [temp_w*3-1:0] v462obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU462 (.l(l[462*data_w +:data_w]), .r(v462ibus), .q(v462obus), .dec(dec[462]));
wire [data_w*3-1:0] v463ibus;
wire [temp_w*3-1:0] v463obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU463 (.l(l[463*data_w +:data_w]), .r(v463ibus), .q(v463obus), .dec(dec[463]));
wire [data_w*3-1:0] v464ibus;
wire [temp_w*3-1:0] v464obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU464 (.l(l[464*data_w +:data_w]), .r(v464ibus), .q(v464obus), .dec(dec[464]));
wire [data_w*3-1:0] v465ibus;
wire [temp_w*3-1:0] v465obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU465 (.l(l[465*data_w +:data_w]), .r(v465ibus), .q(v465obus), .dec(dec[465]));
wire [data_w*3-1:0] v466ibus;
wire [temp_w*3-1:0] v466obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU466 (.l(l[466*data_w +:data_w]), .r(v466ibus), .q(v466obus), .dec(dec[466]));
wire [data_w*3-1:0] v467ibus;
wire [temp_w*3-1:0] v467obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU467 (.l(l[467*data_w +:data_w]), .r(v467ibus), .q(v467obus), .dec(dec[467]));
wire [data_w*3-1:0] v468ibus;
wire [temp_w*3-1:0] v468obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU468 (.l(l[468*data_w +:data_w]), .r(v468ibus), .q(v468obus), .dec(dec[468]));
wire [data_w*3-1:0] v469ibus;
wire [temp_w*3-1:0] v469obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU469 (.l(l[469*data_w +:data_w]), .r(v469ibus), .q(v469obus), .dec(dec[469]));
wire [data_w*3-1:0] v470ibus;
wire [temp_w*3-1:0] v470obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU470 (.l(l[470*data_w +:data_w]), .r(v470ibus), .q(v470obus), .dec(dec[470]));
wire [data_w*3-1:0] v471ibus;
wire [temp_w*3-1:0] v471obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU471 (.l(l[471*data_w +:data_w]), .r(v471ibus), .q(v471obus), .dec(dec[471]));
wire [data_w*3-1:0] v472ibus;
wire [temp_w*3-1:0] v472obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU472 (.l(l[472*data_w +:data_w]), .r(v472ibus), .q(v472obus), .dec(dec[472]));
wire [data_w*3-1:0] v473ibus;
wire [temp_w*3-1:0] v473obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU473 (.l(l[473*data_w +:data_w]), .r(v473ibus), .q(v473obus), .dec(dec[473]));
wire [data_w*3-1:0] v474ibus;
wire [temp_w*3-1:0] v474obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU474 (.l(l[474*data_w +:data_w]), .r(v474ibus), .q(v474obus), .dec(dec[474]));
wire [data_w*3-1:0] v475ibus;
wire [temp_w*3-1:0] v475obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU475 (.l(l[475*data_w +:data_w]), .r(v475ibus), .q(v475obus), .dec(dec[475]));
wire [data_w*3-1:0] v476ibus;
wire [temp_w*3-1:0] v476obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU476 (.l(l[476*data_w +:data_w]), .r(v476ibus), .q(v476obus), .dec(dec[476]));
wire [data_w*3-1:0] v477ibus;
wire [temp_w*3-1:0] v477obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU477 (.l(l[477*data_w +:data_w]), .r(v477ibus), .q(v477obus), .dec(dec[477]));
wire [data_w*3-1:0] v478ibus;
wire [temp_w*3-1:0] v478obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU478 (.l(l[478*data_w +:data_w]), .r(v478ibus), .q(v478obus), .dec(dec[478]));
wire [data_w*3-1:0] v479ibus;
wire [temp_w*3-1:0] v479obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU479 (.l(l[479*data_w +:data_w]), .r(v479ibus), .q(v479obus), .dec(dec[479]));
wire [data_w*6-1:0] v480ibus;
wire [temp_w*6-1:0] v480obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU480 (.l(l[480*data_w +:data_w]), .r(v480ibus), .q(v480obus), .dec(dec[480]));
wire [data_w*6-1:0] v481ibus;
wire [temp_w*6-1:0] v481obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU481 (.l(l[481*data_w +:data_w]), .r(v481ibus), .q(v481obus), .dec(dec[481]));
wire [data_w*6-1:0] v482ibus;
wire [temp_w*6-1:0] v482obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU482 (.l(l[482*data_w +:data_w]), .r(v482ibus), .q(v482obus), .dec(dec[482]));
wire [data_w*6-1:0] v483ibus;
wire [temp_w*6-1:0] v483obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU483 (.l(l[483*data_w +:data_w]), .r(v483ibus), .q(v483obus), .dec(dec[483]));
wire [data_w*6-1:0] v484ibus;
wire [temp_w*6-1:0] v484obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU484 (.l(l[484*data_w +:data_w]), .r(v484ibus), .q(v484obus), .dec(dec[484]));
wire [data_w*6-1:0] v485ibus;
wire [temp_w*6-1:0] v485obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU485 (.l(l[485*data_w +:data_w]), .r(v485ibus), .q(v485obus), .dec(dec[485]));
wire [data_w*6-1:0] v486ibus;
wire [temp_w*6-1:0] v486obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU486 (.l(l[486*data_w +:data_w]), .r(v486ibus), .q(v486obus), .dec(dec[486]));
wire [data_w*6-1:0] v487ibus;
wire [temp_w*6-1:0] v487obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU487 (.l(l[487*data_w +:data_w]), .r(v487ibus), .q(v487obus), .dec(dec[487]));
wire [data_w*6-1:0] v488ibus;
wire [temp_w*6-1:0] v488obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU488 (.l(l[488*data_w +:data_w]), .r(v488ibus), .q(v488obus), .dec(dec[488]));
wire [data_w*6-1:0] v489ibus;
wire [temp_w*6-1:0] v489obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU489 (.l(l[489*data_w +:data_w]), .r(v489ibus), .q(v489obus), .dec(dec[489]));
wire [data_w*6-1:0] v490ibus;
wire [temp_w*6-1:0] v490obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU490 (.l(l[490*data_w +:data_w]), .r(v490ibus), .q(v490obus), .dec(dec[490]));
wire [data_w*6-1:0] v491ibus;
wire [temp_w*6-1:0] v491obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU491 (.l(l[491*data_w +:data_w]), .r(v491ibus), .q(v491obus), .dec(dec[491]));
wire [data_w*6-1:0] v492ibus;
wire [temp_w*6-1:0] v492obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU492 (.l(l[492*data_w +:data_w]), .r(v492ibus), .q(v492obus), .dec(dec[492]));
wire [data_w*6-1:0] v493ibus;
wire [temp_w*6-1:0] v493obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU493 (.l(l[493*data_w +:data_w]), .r(v493ibus), .q(v493obus), .dec(dec[493]));
wire [data_w*6-1:0] v494ibus;
wire [temp_w*6-1:0] v494obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU494 (.l(l[494*data_w +:data_w]), .r(v494ibus), .q(v494obus), .dec(dec[494]));
wire [data_w*6-1:0] v495ibus;
wire [temp_w*6-1:0] v495obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU495 (.l(l[495*data_w +:data_w]), .r(v495ibus), .q(v495obus), .dec(dec[495]));
wire [data_w*6-1:0] v496ibus;
wire [temp_w*6-1:0] v496obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU496 (.l(l[496*data_w +:data_w]), .r(v496ibus), .q(v496obus), .dec(dec[496]));
wire [data_w*6-1:0] v497ibus;
wire [temp_w*6-1:0] v497obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU497 (.l(l[497*data_w +:data_w]), .r(v497ibus), .q(v497obus), .dec(dec[497]));
wire [data_w*6-1:0] v498ibus;
wire [temp_w*6-1:0] v498obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU498 (.l(l[498*data_w +:data_w]), .r(v498ibus), .q(v498obus), .dec(dec[498]));
wire [data_w*6-1:0] v499ibus;
wire [temp_w*6-1:0] v499obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU499 (.l(l[499*data_w +:data_w]), .r(v499ibus), .q(v499obus), .dec(dec[499]));
wire [data_w*6-1:0] v500ibus;
wire [temp_w*6-1:0] v500obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU500 (.l(l[500*data_w +:data_w]), .r(v500ibus), .q(v500obus), .dec(dec[500]));
wire [data_w*6-1:0] v501ibus;
wire [temp_w*6-1:0] v501obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU501 (.l(l[501*data_w +:data_w]), .r(v501ibus), .q(v501obus), .dec(dec[501]));
wire [data_w*6-1:0] v502ibus;
wire [temp_w*6-1:0] v502obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU502 (.l(l[502*data_w +:data_w]), .r(v502ibus), .q(v502obus), .dec(dec[502]));
wire [data_w*6-1:0] v503ibus;
wire [temp_w*6-1:0] v503obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU503 (.l(l[503*data_w +:data_w]), .r(v503ibus), .q(v503obus), .dec(dec[503]));
wire [data_w*6-1:0] v504ibus;
wire [temp_w*6-1:0] v504obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU504 (.l(l[504*data_w +:data_w]), .r(v504ibus), .q(v504obus), .dec(dec[504]));
wire [data_w*6-1:0] v505ibus;
wire [temp_w*6-1:0] v505obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU505 (.l(l[505*data_w +:data_w]), .r(v505ibus), .q(v505obus), .dec(dec[505]));
wire [data_w*6-1:0] v506ibus;
wire [temp_w*6-1:0] v506obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU506 (.l(l[506*data_w +:data_w]), .r(v506ibus), .q(v506obus), .dec(dec[506]));
wire [data_w*6-1:0] v507ibus;
wire [temp_w*6-1:0] v507obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU507 (.l(l[507*data_w +:data_w]), .r(v507ibus), .q(v507obus), .dec(dec[507]));
wire [data_w*6-1:0] v508ibus;
wire [temp_w*6-1:0] v508obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU508 (.l(l[508*data_w +:data_w]), .r(v508ibus), .q(v508obus), .dec(dec[508]));
wire [data_w*6-1:0] v509ibus;
wire [temp_w*6-1:0] v509obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU509 (.l(l[509*data_w +:data_w]), .r(v509ibus), .q(v509obus), .dec(dec[509]));
wire [data_w*6-1:0] v510ibus;
wire [temp_w*6-1:0] v510obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU510 (.l(l[510*data_w +:data_w]), .r(v510ibus), .q(v510obus), .dec(dec[510]));
wire [data_w*6-1:0] v511ibus;
wire [temp_w*6-1:0] v511obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU511 (.l(l[511*data_w +:data_w]), .r(v511ibus), .q(v511obus), .dec(dec[511]));
wire [data_w*6-1:0] v512ibus;
wire [temp_w*6-1:0] v512obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU512 (.l(l[512*data_w +:data_w]), .r(v512ibus), .q(v512obus), .dec(dec[512]));
wire [data_w*6-1:0] v513ibus;
wire [temp_w*6-1:0] v513obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU513 (.l(l[513*data_w +:data_w]), .r(v513ibus), .q(v513obus), .dec(dec[513]));
wire [data_w*6-1:0] v514ibus;
wire [temp_w*6-1:0] v514obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU514 (.l(l[514*data_w +:data_w]), .r(v514ibus), .q(v514obus), .dec(dec[514]));
wire [data_w*6-1:0] v515ibus;
wire [temp_w*6-1:0] v515obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU515 (.l(l[515*data_w +:data_w]), .r(v515ibus), .q(v515obus), .dec(dec[515]));
wire [data_w*6-1:0] v516ibus;
wire [temp_w*6-1:0] v516obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU516 (.l(l[516*data_w +:data_w]), .r(v516ibus), .q(v516obus), .dec(dec[516]));
wire [data_w*6-1:0] v517ibus;
wire [temp_w*6-1:0] v517obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU517 (.l(l[517*data_w +:data_w]), .r(v517ibus), .q(v517obus), .dec(dec[517]));
wire [data_w*6-1:0] v518ibus;
wire [temp_w*6-1:0] v518obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU518 (.l(l[518*data_w +:data_w]), .r(v518ibus), .q(v518obus), .dec(dec[518]));
wire [data_w*6-1:0] v519ibus;
wire [temp_w*6-1:0] v519obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU519 (.l(l[519*data_w +:data_w]), .r(v519ibus), .q(v519obus), .dec(dec[519]));
wire [data_w*6-1:0] v520ibus;
wire [temp_w*6-1:0] v520obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU520 (.l(l[520*data_w +:data_w]), .r(v520ibus), .q(v520obus), .dec(dec[520]));
wire [data_w*6-1:0] v521ibus;
wire [temp_w*6-1:0] v521obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU521 (.l(l[521*data_w +:data_w]), .r(v521ibus), .q(v521obus), .dec(dec[521]));
wire [data_w*6-1:0] v522ibus;
wire [temp_w*6-1:0] v522obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU522 (.l(l[522*data_w +:data_w]), .r(v522ibus), .q(v522obus), .dec(dec[522]));
wire [data_w*6-1:0] v523ibus;
wire [temp_w*6-1:0] v523obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU523 (.l(l[523*data_w +:data_w]), .r(v523ibus), .q(v523obus), .dec(dec[523]));
wire [data_w*6-1:0] v524ibus;
wire [temp_w*6-1:0] v524obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU524 (.l(l[524*data_w +:data_w]), .r(v524ibus), .q(v524obus), .dec(dec[524]));
wire [data_w*6-1:0] v525ibus;
wire [temp_w*6-1:0] v525obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU525 (.l(l[525*data_w +:data_w]), .r(v525ibus), .q(v525obus), .dec(dec[525]));
wire [data_w*6-1:0] v526ibus;
wire [temp_w*6-1:0] v526obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU526 (.l(l[526*data_w +:data_w]), .r(v526ibus), .q(v526obus), .dec(dec[526]));
wire [data_w*6-1:0] v527ibus;
wire [temp_w*6-1:0] v527obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU527 (.l(l[527*data_w +:data_w]), .r(v527ibus), .q(v527obus), .dec(dec[527]));
wire [data_w*6-1:0] v528ibus;
wire [temp_w*6-1:0] v528obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU528 (.l(l[528*data_w +:data_w]), .r(v528ibus), .q(v528obus), .dec(dec[528]));
wire [data_w*6-1:0] v529ibus;
wire [temp_w*6-1:0] v529obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU529 (.l(l[529*data_w +:data_w]), .r(v529ibus), .q(v529obus), .dec(dec[529]));
wire [data_w*6-1:0] v530ibus;
wire [temp_w*6-1:0] v530obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU530 (.l(l[530*data_w +:data_w]), .r(v530ibus), .q(v530obus), .dec(dec[530]));
wire [data_w*6-1:0] v531ibus;
wire [temp_w*6-1:0] v531obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU531 (.l(l[531*data_w +:data_w]), .r(v531ibus), .q(v531obus), .dec(dec[531]));
wire [data_w*6-1:0] v532ibus;
wire [temp_w*6-1:0] v532obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU532 (.l(l[532*data_w +:data_w]), .r(v532ibus), .q(v532obus), .dec(dec[532]));
wire [data_w*6-1:0] v533ibus;
wire [temp_w*6-1:0] v533obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU533 (.l(l[533*data_w +:data_w]), .r(v533ibus), .q(v533obus), .dec(dec[533]));
wire [data_w*6-1:0] v534ibus;
wire [temp_w*6-1:0] v534obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU534 (.l(l[534*data_w +:data_w]), .r(v534ibus), .q(v534obus), .dec(dec[534]));
wire [data_w*6-1:0] v535ibus;
wire [temp_w*6-1:0] v535obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU535 (.l(l[535*data_w +:data_w]), .r(v535ibus), .q(v535obus), .dec(dec[535]));
wire [data_w*6-1:0] v536ibus;
wire [temp_w*6-1:0] v536obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU536 (.l(l[536*data_w +:data_w]), .r(v536ibus), .q(v536obus), .dec(dec[536]));
wire [data_w*6-1:0] v537ibus;
wire [temp_w*6-1:0] v537obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU537 (.l(l[537*data_w +:data_w]), .r(v537ibus), .q(v537obus), .dec(dec[537]));
wire [data_w*6-1:0] v538ibus;
wire [temp_w*6-1:0] v538obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU538 (.l(l[538*data_w +:data_w]), .r(v538ibus), .q(v538obus), .dec(dec[538]));
wire [data_w*6-1:0] v539ibus;
wire [temp_w*6-1:0] v539obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU539 (.l(l[539*data_w +:data_w]), .r(v539ibus), .q(v539obus), .dec(dec[539]));
wire [data_w*6-1:0] v540ibus;
wire [temp_w*6-1:0] v540obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU540 (.l(l[540*data_w +:data_w]), .r(v540ibus), .q(v540obus), .dec(dec[540]));
wire [data_w*6-1:0] v541ibus;
wire [temp_w*6-1:0] v541obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU541 (.l(l[541*data_w +:data_w]), .r(v541ibus), .q(v541obus), .dec(dec[541]));
wire [data_w*6-1:0] v542ibus;
wire [temp_w*6-1:0] v542obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU542 (.l(l[542*data_w +:data_w]), .r(v542ibus), .q(v542obus), .dec(dec[542]));
wire [data_w*6-1:0] v543ibus;
wire [temp_w*6-1:0] v543obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU543 (.l(l[543*data_w +:data_w]), .r(v543ibus), .q(v543obus), .dec(dec[543]));
wire [data_w*6-1:0] v544ibus;
wire [temp_w*6-1:0] v544obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU544 (.l(l[544*data_w +:data_w]), .r(v544ibus), .q(v544obus), .dec(dec[544]));
wire [data_w*6-1:0] v545ibus;
wire [temp_w*6-1:0] v545obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU545 (.l(l[545*data_w +:data_w]), .r(v545ibus), .q(v545obus), .dec(dec[545]));
wire [data_w*6-1:0] v546ibus;
wire [temp_w*6-1:0] v546obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU546 (.l(l[546*data_w +:data_w]), .r(v546ibus), .q(v546obus), .dec(dec[546]));
wire [data_w*6-1:0] v547ibus;
wire [temp_w*6-1:0] v547obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU547 (.l(l[547*data_w +:data_w]), .r(v547ibus), .q(v547obus), .dec(dec[547]));
wire [data_w*6-1:0] v548ibus;
wire [temp_w*6-1:0] v548obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU548 (.l(l[548*data_w +:data_w]), .r(v548ibus), .q(v548obus), .dec(dec[548]));
wire [data_w*6-1:0] v549ibus;
wire [temp_w*6-1:0] v549obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU549 (.l(l[549*data_w +:data_w]), .r(v549ibus), .q(v549obus), .dec(dec[549]));
wire [data_w*6-1:0] v550ibus;
wire [temp_w*6-1:0] v550obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU550 (.l(l[550*data_w +:data_w]), .r(v550ibus), .q(v550obus), .dec(dec[550]));
wire [data_w*6-1:0] v551ibus;
wire [temp_w*6-1:0] v551obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU551 (.l(l[551*data_w +:data_w]), .r(v551ibus), .q(v551obus), .dec(dec[551]));
wire [data_w*6-1:0] v552ibus;
wire [temp_w*6-1:0] v552obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU552 (.l(l[552*data_w +:data_w]), .r(v552ibus), .q(v552obus), .dec(dec[552]));
wire [data_w*6-1:0] v553ibus;
wire [temp_w*6-1:0] v553obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU553 (.l(l[553*data_w +:data_w]), .r(v553ibus), .q(v553obus), .dec(dec[553]));
wire [data_w*6-1:0] v554ibus;
wire [temp_w*6-1:0] v554obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU554 (.l(l[554*data_w +:data_w]), .r(v554ibus), .q(v554obus), .dec(dec[554]));
wire [data_w*6-1:0] v555ibus;
wire [temp_w*6-1:0] v555obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU555 (.l(l[555*data_w +:data_w]), .r(v555ibus), .q(v555obus), .dec(dec[555]));
wire [data_w*6-1:0] v556ibus;
wire [temp_w*6-1:0] v556obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU556 (.l(l[556*data_w +:data_w]), .r(v556ibus), .q(v556obus), .dec(dec[556]));
wire [data_w*6-1:0] v557ibus;
wire [temp_w*6-1:0] v557obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU557 (.l(l[557*data_w +:data_w]), .r(v557ibus), .q(v557obus), .dec(dec[557]));
wire [data_w*6-1:0] v558ibus;
wire [temp_w*6-1:0] v558obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU558 (.l(l[558*data_w +:data_w]), .r(v558ibus), .q(v558obus), .dec(dec[558]));
wire [data_w*6-1:0] v559ibus;
wire [temp_w*6-1:0] v559obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU559 (.l(l[559*data_w +:data_w]), .r(v559ibus), .q(v559obus), .dec(dec[559]));
wire [data_w*6-1:0] v560ibus;
wire [temp_w*6-1:0] v560obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU560 (.l(l[560*data_w +:data_w]), .r(v560ibus), .q(v560obus), .dec(dec[560]));
wire [data_w*6-1:0] v561ibus;
wire [temp_w*6-1:0] v561obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU561 (.l(l[561*data_w +:data_w]), .r(v561ibus), .q(v561obus), .dec(dec[561]));
wire [data_w*6-1:0] v562ibus;
wire [temp_w*6-1:0] v562obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU562 (.l(l[562*data_w +:data_w]), .r(v562ibus), .q(v562obus), .dec(dec[562]));
wire [data_w*6-1:0] v563ibus;
wire [temp_w*6-1:0] v563obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU563 (.l(l[563*data_w +:data_w]), .r(v563ibus), .q(v563obus), .dec(dec[563]));
wire [data_w*6-1:0] v564ibus;
wire [temp_w*6-1:0] v564obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU564 (.l(l[564*data_w +:data_w]), .r(v564ibus), .q(v564obus), .dec(dec[564]));
wire [data_w*6-1:0] v565ibus;
wire [temp_w*6-1:0] v565obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU565 (.l(l[565*data_w +:data_w]), .r(v565ibus), .q(v565obus), .dec(dec[565]));
wire [data_w*6-1:0] v566ibus;
wire [temp_w*6-1:0] v566obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU566 (.l(l[566*data_w +:data_w]), .r(v566ibus), .q(v566obus), .dec(dec[566]));
wire [data_w*6-1:0] v567ibus;
wire [temp_w*6-1:0] v567obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU567 (.l(l[567*data_w +:data_w]), .r(v567ibus), .q(v567obus), .dec(dec[567]));
wire [data_w*6-1:0] v568ibus;
wire [temp_w*6-1:0] v568obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU568 (.l(l[568*data_w +:data_w]), .r(v568ibus), .q(v568obus), .dec(dec[568]));
wire [data_w*6-1:0] v569ibus;
wire [temp_w*6-1:0] v569obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU569 (.l(l[569*data_w +:data_w]), .r(v569ibus), .q(v569obus), .dec(dec[569]));
wire [data_w*6-1:0] v570ibus;
wire [temp_w*6-1:0] v570obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU570 (.l(l[570*data_w +:data_w]), .r(v570ibus), .q(v570obus), .dec(dec[570]));
wire [data_w*6-1:0] v571ibus;
wire [temp_w*6-1:0] v571obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU571 (.l(l[571*data_w +:data_w]), .r(v571ibus), .q(v571obus), .dec(dec[571]));
wire [data_w*6-1:0] v572ibus;
wire [temp_w*6-1:0] v572obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU572 (.l(l[572*data_w +:data_w]), .r(v572ibus), .q(v572obus), .dec(dec[572]));
wire [data_w*6-1:0] v573ibus;
wire [temp_w*6-1:0] v573obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU573 (.l(l[573*data_w +:data_w]), .r(v573ibus), .q(v573obus), .dec(dec[573]));
wire [data_w*6-1:0] v574ibus;
wire [temp_w*6-1:0] v574obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU574 (.l(l[574*data_w +:data_w]), .r(v574ibus), .q(v574obus), .dec(dec[574]));
wire [data_w*6-1:0] v575ibus;
wire [temp_w*6-1:0] v575obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU575 (.l(l[575*data_w +:data_w]), .r(v575ibus), .q(v575obus), .dec(dec[575]));
wire [data_w*3-1:0] v576ibus;
wire [temp_w*3-1:0] v576obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU576 (.l(l[576*data_w +:data_w]), .r(v576ibus), .q(v576obus), .dec(dec[576]));
wire [data_w*3-1:0] v577ibus;
wire [temp_w*3-1:0] v577obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU577 (.l(l[577*data_w +:data_w]), .r(v577ibus), .q(v577obus), .dec(dec[577]));
wire [data_w*3-1:0] v578ibus;
wire [temp_w*3-1:0] v578obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU578 (.l(l[578*data_w +:data_w]), .r(v578ibus), .q(v578obus), .dec(dec[578]));
wire [data_w*3-1:0] v579ibus;
wire [temp_w*3-1:0] v579obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU579 (.l(l[579*data_w +:data_w]), .r(v579ibus), .q(v579obus), .dec(dec[579]));
wire [data_w*3-1:0] v580ibus;
wire [temp_w*3-1:0] v580obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU580 (.l(l[580*data_w +:data_w]), .r(v580ibus), .q(v580obus), .dec(dec[580]));
wire [data_w*3-1:0] v581ibus;
wire [temp_w*3-1:0] v581obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU581 (.l(l[581*data_w +:data_w]), .r(v581ibus), .q(v581obus), .dec(dec[581]));
wire [data_w*3-1:0] v582ibus;
wire [temp_w*3-1:0] v582obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU582 (.l(l[582*data_w +:data_w]), .r(v582ibus), .q(v582obus), .dec(dec[582]));
wire [data_w*3-1:0] v583ibus;
wire [temp_w*3-1:0] v583obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU583 (.l(l[583*data_w +:data_w]), .r(v583ibus), .q(v583obus), .dec(dec[583]));
wire [data_w*3-1:0] v584ibus;
wire [temp_w*3-1:0] v584obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU584 (.l(l[584*data_w +:data_w]), .r(v584ibus), .q(v584obus), .dec(dec[584]));
wire [data_w*3-1:0] v585ibus;
wire [temp_w*3-1:0] v585obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU585 (.l(l[585*data_w +:data_w]), .r(v585ibus), .q(v585obus), .dec(dec[585]));
wire [data_w*3-1:0] v586ibus;
wire [temp_w*3-1:0] v586obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU586 (.l(l[586*data_w +:data_w]), .r(v586ibus), .q(v586obus), .dec(dec[586]));
wire [data_w*3-1:0] v587ibus;
wire [temp_w*3-1:0] v587obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU587 (.l(l[587*data_w +:data_w]), .r(v587ibus), .q(v587obus), .dec(dec[587]));
wire [data_w*3-1:0] v588ibus;
wire [temp_w*3-1:0] v588obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU588 (.l(l[588*data_w +:data_w]), .r(v588ibus), .q(v588obus), .dec(dec[588]));
wire [data_w*3-1:0] v589ibus;
wire [temp_w*3-1:0] v589obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU589 (.l(l[589*data_w +:data_w]), .r(v589ibus), .q(v589obus), .dec(dec[589]));
wire [data_w*3-1:0] v590ibus;
wire [temp_w*3-1:0] v590obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU590 (.l(l[590*data_w +:data_w]), .r(v590ibus), .q(v590obus), .dec(dec[590]));
wire [data_w*3-1:0] v591ibus;
wire [temp_w*3-1:0] v591obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU591 (.l(l[591*data_w +:data_w]), .r(v591ibus), .q(v591obus), .dec(dec[591]));
wire [data_w*3-1:0] v592ibus;
wire [temp_w*3-1:0] v592obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU592 (.l(l[592*data_w +:data_w]), .r(v592ibus), .q(v592obus), .dec(dec[592]));
wire [data_w*3-1:0] v593ibus;
wire [temp_w*3-1:0] v593obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU593 (.l(l[593*data_w +:data_w]), .r(v593ibus), .q(v593obus), .dec(dec[593]));
wire [data_w*3-1:0] v594ibus;
wire [temp_w*3-1:0] v594obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU594 (.l(l[594*data_w +:data_w]), .r(v594ibus), .q(v594obus), .dec(dec[594]));
wire [data_w*3-1:0] v595ibus;
wire [temp_w*3-1:0] v595obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU595 (.l(l[595*data_w +:data_w]), .r(v595ibus), .q(v595obus), .dec(dec[595]));
wire [data_w*3-1:0] v596ibus;
wire [temp_w*3-1:0] v596obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU596 (.l(l[596*data_w +:data_w]), .r(v596ibus), .q(v596obus), .dec(dec[596]));
wire [data_w*3-1:0] v597ibus;
wire [temp_w*3-1:0] v597obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU597 (.l(l[597*data_w +:data_w]), .r(v597ibus), .q(v597obus), .dec(dec[597]));
wire [data_w*3-1:0] v598ibus;
wire [temp_w*3-1:0] v598obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU598 (.l(l[598*data_w +:data_w]), .r(v598ibus), .q(v598obus), .dec(dec[598]));
wire [data_w*3-1:0] v599ibus;
wire [temp_w*3-1:0] v599obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU599 (.l(l[599*data_w +:data_w]), .r(v599ibus), .q(v599obus), .dec(dec[599]));
wire [data_w*3-1:0] v600ibus;
wire [temp_w*3-1:0] v600obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU600 (.l(l[600*data_w +:data_w]), .r(v600ibus), .q(v600obus), .dec(dec[600]));
wire [data_w*3-1:0] v601ibus;
wire [temp_w*3-1:0] v601obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU601 (.l(l[601*data_w +:data_w]), .r(v601ibus), .q(v601obus), .dec(dec[601]));
wire [data_w*3-1:0] v602ibus;
wire [temp_w*3-1:0] v602obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU602 (.l(l[602*data_w +:data_w]), .r(v602ibus), .q(v602obus), .dec(dec[602]));
wire [data_w*3-1:0] v603ibus;
wire [temp_w*3-1:0] v603obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU603 (.l(l[603*data_w +:data_w]), .r(v603ibus), .q(v603obus), .dec(dec[603]));
wire [data_w*3-1:0] v604ibus;
wire [temp_w*3-1:0] v604obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU604 (.l(l[604*data_w +:data_w]), .r(v604ibus), .q(v604obus), .dec(dec[604]));
wire [data_w*3-1:0] v605ibus;
wire [temp_w*3-1:0] v605obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU605 (.l(l[605*data_w +:data_w]), .r(v605ibus), .q(v605obus), .dec(dec[605]));
wire [data_w*3-1:0] v606ibus;
wire [temp_w*3-1:0] v606obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU606 (.l(l[606*data_w +:data_w]), .r(v606ibus), .q(v606obus), .dec(dec[606]));
wire [data_w*3-1:0] v607ibus;
wire [temp_w*3-1:0] v607obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU607 (.l(l[607*data_w +:data_w]), .r(v607ibus), .q(v607obus), .dec(dec[607]));
wire [data_w*3-1:0] v608ibus;
wire [temp_w*3-1:0] v608obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU608 (.l(l[608*data_w +:data_w]), .r(v608ibus), .q(v608obus), .dec(dec[608]));
wire [data_w*3-1:0] v609ibus;
wire [temp_w*3-1:0] v609obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU609 (.l(l[609*data_w +:data_w]), .r(v609ibus), .q(v609obus), .dec(dec[609]));
wire [data_w*3-1:0] v610ibus;
wire [temp_w*3-1:0] v610obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU610 (.l(l[610*data_w +:data_w]), .r(v610ibus), .q(v610obus), .dec(dec[610]));
wire [data_w*3-1:0] v611ibus;
wire [temp_w*3-1:0] v611obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU611 (.l(l[611*data_w +:data_w]), .r(v611ibus), .q(v611obus), .dec(dec[611]));
wire [data_w*3-1:0] v612ibus;
wire [temp_w*3-1:0] v612obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU612 (.l(l[612*data_w +:data_w]), .r(v612ibus), .q(v612obus), .dec(dec[612]));
wire [data_w*3-1:0] v613ibus;
wire [temp_w*3-1:0] v613obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU613 (.l(l[613*data_w +:data_w]), .r(v613ibus), .q(v613obus), .dec(dec[613]));
wire [data_w*3-1:0] v614ibus;
wire [temp_w*3-1:0] v614obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU614 (.l(l[614*data_w +:data_w]), .r(v614ibus), .q(v614obus), .dec(dec[614]));
wire [data_w*3-1:0] v615ibus;
wire [temp_w*3-1:0] v615obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU615 (.l(l[615*data_w +:data_w]), .r(v615ibus), .q(v615obus), .dec(dec[615]));
wire [data_w*3-1:0] v616ibus;
wire [temp_w*3-1:0] v616obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU616 (.l(l[616*data_w +:data_w]), .r(v616ibus), .q(v616obus), .dec(dec[616]));
wire [data_w*3-1:0] v617ibus;
wire [temp_w*3-1:0] v617obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU617 (.l(l[617*data_w +:data_w]), .r(v617ibus), .q(v617obus), .dec(dec[617]));
wire [data_w*3-1:0] v618ibus;
wire [temp_w*3-1:0] v618obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU618 (.l(l[618*data_w +:data_w]), .r(v618ibus), .q(v618obus), .dec(dec[618]));
wire [data_w*3-1:0] v619ibus;
wire [temp_w*3-1:0] v619obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU619 (.l(l[619*data_w +:data_w]), .r(v619ibus), .q(v619obus), .dec(dec[619]));
wire [data_w*3-1:0] v620ibus;
wire [temp_w*3-1:0] v620obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU620 (.l(l[620*data_w +:data_w]), .r(v620ibus), .q(v620obus), .dec(dec[620]));
wire [data_w*3-1:0] v621ibus;
wire [temp_w*3-1:0] v621obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU621 (.l(l[621*data_w +:data_w]), .r(v621ibus), .q(v621obus), .dec(dec[621]));
wire [data_w*3-1:0] v622ibus;
wire [temp_w*3-1:0] v622obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU622 (.l(l[622*data_w +:data_w]), .r(v622ibus), .q(v622obus), .dec(dec[622]));
wire [data_w*3-1:0] v623ibus;
wire [temp_w*3-1:0] v623obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU623 (.l(l[623*data_w +:data_w]), .r(v623ibus), .q(v623obus), .dec(dec[623]));
wire [data_w*3-1:0] v624ibus;
wire [temp_w*3-1:0] v624obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU624 (.l(l[624*data_w +:data_w]), .r(v624ibus), .q(v624obus), .dec(dec[624]));
wire [data_w*3-1:0] v625ibus;
wire [temp_w*3-1:0] v625obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU625 (.l(l[625*data_w +:data_w]), .r(v625ibus), .q(v625obus), .dec(dec[625]));
wire [data_w*3-1:0] v626ibus;
wire [temp_w*3-1:0] v626obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU626 (.l(l[626*data_w +:data_w]), .r(v626ibus), .q(v626obus), .dec(dec[626]));
wire [data_w*3-1:0] v627ibus;
wire [temp_w*3-1:0] v627obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU627 (.l(l[627*data_w +:data_w]), .r(v627ibus), .q(v627obus), .dec(dec[627]));
wire [data_w*3-1:0] v628ibus;
wire [temp_w*3-1:0] v628obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU628 (.l(l[628*data_w +:data_w]), .r(v628ibus), .q(v628obus), .dec(dec[628]));
wire [data_w*3-1:0] v629ibus;
wire [temp_w*3-1:0] v629obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU629 (.l(l[629*data_w +:data_w]), .r(v629ibus), .q(v629obus), .dec(dec[629]));
wire [data_w*3-1:0] v630ibus;
wire [temp_w*3-1:0] v630obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU630 (.l(l[630*data_w +:data_w]), .r(v630ibus), .q(v630obus), .dec(dec[630]));
wire [data_w*3-1:0] v631ibus;
wire [temp_w*3-1:0] v631obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU631 (.l(l[631*data_w +:data_w]), .r(v631ibus), .q(v631obus), .dec(dec[631]));
wire [data_w*3-1:0] v632ibus;
wire [temp_w*3-1:0] v632obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU632 (.l(l[632*data_w +:data_w]), .r(v632ibus), .q(v632obus), .dec(dec[632]));
wire [data_w*3-1:0] v633ibus;
wire [temp_w*3-1:0] v633obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU633 (.l(l[633*data_w +:data_w]), .r(v633ibus), .q(v633obus), .dec(dec[633]));
wire [data_w*3-1:0] v634ibus;
wire [temp_w*3-1:0] v634obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU634 (.l(l[634*data_w +:data_w]), .r(v634ibus), .q(v634obus), .dec(dec[634]));
wire [data_w*3-1:0] v635ibus;
wire [temp_w*3-1:0] v635obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU635 (.l(l[635*data_w +:data_w]), .r(v635ibus), .q(v635obus), .dec(dec[635]));
wire [data_w*3-1:0] v636ibus;
wire [temp_w*3-1:0] v636obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU636 (.l(l[636*data_w +:data_w]), .r(v636ibus), .q(v636obus), .dec(dec[636]));
wire [data_w*3-1:0] v637ibus;
wire [temp_w*3-1:0] v637obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU637 (.l(l[637*data_w +:data_w]), .r(v637ibus), .q(v637obus), .dec(dec[637]));
wire [data_w*3-1:0] v638ibus;
wire [temp_w*3-1:0] v638obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU638 (.l(l[638*data_w +:data_w]), .r(v638ibus), .q(v638obus), .dec(dec[638]));
wire [data_w*3-1:0] v639ibus;
wire [temp_w*3-1:0] v639obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU639 (.l(l[639*data_w +:data_w]), .r(v639ibus), .q(v639obus), .dec(dec[639]));
wire [data_w*3-1:0] v640ibus;
wire [temp_w*3-1:0] v640obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU640 (.l(l[640*data_w +:data_w]), .r(v640ibus), .q(v640obus), .dec(dec[640]));
wire [data_w*3-1:0] v641ibus;
wire [temp_w*3-1:0] v641obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU641 (.l(l[641*data_w +:data_w]), .r(v641ibus), .q(v641obus), .dec(dec[641]));
wire [data_w*3-1:0] v642ibus;
wire [temp_w*3-1:0] v642obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU642 (.l(l[642*data_w +:data_w]), .r(v642ibus), .q(v642obus), .dec(dec[642]));
wire [data_w*3-1:0] v643ibus;
wire [temp_w*3-1:0] v643obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU643 (.l(l[643*data_w +:data_w]), .r(v643ibus), .q(v643obus), .dec(dec[643]));
wire [data_w*3-1:0] v644ibus;
wire [temp_w*3-1:0] v644obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU644 (.l(l[644*data_w +:data_w]), .r(v644ibus), .q(v644obus), .dec(dec[644]));
wire [data_w*3-1:0] v645ibus;
wire [temp_w*3-1:0] v645obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU645 (.l(l[645*data_w +:data_w]), .r(v645ibus), .q(v645obus), .dec(dec[645]));
wire [data_w*3-1:0] v646ibus;
wire [temp_w*3-1:0] v646obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU646 (.l(l[646*data_w +:data_w]), .r(v646ibus), .q(v646obus), .dec(dec[646]));
wire [data_w*3-1:0] v647ibus;
wire [temp_w*3-1:0] v647obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU647 (.l(l[647*data_w +:data_w]), .r(v647ibus), .q(v647obus), .dec(dec[647]));
wire [data_w*3-1:0] v648ibus;
wire [temp_w*3-1:0] v648obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU648 (.l(l[648*data_w +:data_w]), .r(v648ibus), .q(v648obus), .dec(dec[648]));
wire [data_w*3-1:0] v649ibus;
wire [temp_w*3-1:0] v649obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU649 (.l(l[649*data_w +:data_w]), .r(v649ibus), .q(v649obus), .dec(dec[649]));
wire [data_w*3-1:0] v650ibus;
wire [temp_w*3-1:0] v650obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU650 (.l(l[650*data_w +:data_w]), .r(v650ibus), .q(v650obus), .dec(dec[650]));
wire [data_w*3-1:0] v651ibus;
wire [temp_w*3-1:0] v651obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU651 (.l(l[651*data_w +:data_w]), .r(v651ibus), .q(v651obus), .dec(dec[651]));
wire [data_w*3-1:0] v652ibus;
wire [temp_w*3-1:0] v652obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU652 (.l(l[652*data_w +:data_w]), .r(v652ibus), .q(v652obus), .dec(dec[652]));
wire [data_w*3-1:0] v653ibus;
wire [temp_w*3-1:0] v653obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU653 (.l(l[653*data_w +:data_w]), .r(v653ibus), .q(v653obus), .dec(dec[653]));
wire [data_w*3-1:0] v654ibus;
wire [temp_w*3-1:0] v654obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU654 (.l(l[654*data_w +:data_w]), .r(v654ibus), .q(v654obus), .dec(dec[654]));
wire [data_w*3-1:0] v655ibus;
wire [temp_w*3-1:0] v655obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU655 (.l(l[655*data_w +:data_w]), .r(v655ibus), .q(v655obus), .dec(dec[655]));
wire [data_w*3-1:0] v656ibus;
wire [temp_w*3-1:0] v656obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU656 (.l(l[656*data_w +:data_w]), .r(v656ibus), .q(v656obus), .dec(dec[656]));
wire [data_w*3-1:0] v657ibus;
wire [temp_w*3-1:0] v657obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU657 (.l(l[657*data_w +:data_w]), .r(v657ibus), .q(v657obus), .dec(dec[657]));
wire [data_w*3-1:0] v658ibus;
wire [temp_w*3-1:0] v658obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU658 (.l(l[658*data_w +:data_w]), .r(v658ibus), .q(v658obus), .dec(dec[658]));
wire [data_w*3-1:0] v659ibus;
wire [temp_w*3-1:0] v659obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU659 (.l(l[659*data_w +:data_w]), .r(v659ibus), .q(v659obus), .dec(dec[659]));
wire [data_w*3-1:0] v660ibus;
wire [temp_w*3-1:0] v660obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU660 (.l(l[660*data_w +:data_w]), .r(v660ibus), .q(v660obus), .dec(dec[660]));
wire [data_w*3-1:0] v661ibus;
wire [temp_w*3-1:0] v661obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU661 (.l(l[661*data_w +:data_w]), .r(v661ibus), .q(v661obus), .dec(dec[661]));
wire [data_w*3-1:0] v662ibus;
wire [temp_w*3-1:0] v662obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU662 (.l(l[662*data_w +:data_w]), .r(v662ibus), .q(v662obus), .dec(dec[662]));
wire [data_w*3-1:0] v663ibus;
wire [temp_w*3-1:0] v663obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU663 (.l(l[663*data_w +:data_w]), .r(v663ibus), .q(v663obus), .dec(dec[663]));
wire [data_w*3-1:0] v664ibus;
wire [temp_w*3-1:0] v664obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU664 (.l(l[664*data_w +:data_w]), .r(v664ibus), .q(v664obus), .dec(dec[664]));
wire [data_w*3-1:0] v665ibus;
wire [temp_w*3-1:0] v665obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU665 (.l(l[665*data_w +:data_w]), .r(v665ibus), .q(v665obus), .dec(dec[665]));
wire [data_w*3-1:0] v666ibus;
wire [temp_w*3-1:0] v666obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU666 (.l(l[666*data_w +:data_w]), .r(v666ibus), .q(v666obus), .dec(dec[666]));
wire [data_w*3-1:0] v667ibus;
wire [temp_w*3-1:0] v667obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU667 (.l(l[667*data_w +:data_w]), .r(v667ibus), .q(v667obus), .dec(dec[667]));
wire [data_w*3-1:0] v668ibus;
wire [temp_w*3-1:0] v668obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU668 (.l(l[668*data_w +:data_w]), .r(v668ibus), .q(v668obus), .dec(dec[668]));
wire [data_w*3-1:0] v669ibus;
wire [temp_w*3-1:0] v669obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU669 (.l(l[669*data_w +:data_w]), .r(v669ibus), .q(v669obus), .dec(dec[669]));
wire [data_w*3-1:0] v670ibus;
wire [temp_w*3-1:0] v670obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU670 (.l(l[670*data_w +:data_w]), .r(v670ibus), .q(v670obus), .dec(dec[670]));
wire [data_w*3-1:0] v671ibus;
wire [temp_w*3-1:0] v671obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU671 (.l(l[671*data_w +:data_w]), .r(v671ibus), .q(v671obus), .dec(dec[671]));
wire [data_w*6-1:0] v672ibus;
wire [temp_w*6-1:0] v672obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU672 (.l(l[672*data_w +:data_w]), .r(v672ibus), .q(v672obus), .dec(dec[672]));
wire [data_w*6-1:0] v673ibus;
wire [temp_w*6-1:0] v673obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU673 (.l(l[673*data_w +:data_w]), .r(v673ibus), .q(v673obus), .dec(dec[673]));
wire [data_w*6-1:0] v674ibus;
wire [temp_w*6-1:0] v674obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU674 (.l(l[674*data_w +:data_w]), .r(v674ibus), .q(v674obus), .dec(dec[674]));
wire [data_w*6-1:0] v675ibus;
wire [temp_w*6-1:0] v675obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU675 (.l(l[675*data_w +:data_w]), .r(v675ibus), .q(v675obus), .dec(dec[675]));
wire [data_w*6-1:0] v676ibus;
wire [temp_w*6-1:0] v676obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU676 (.l(l[676*data_w +:data_w]), .r(v676ibus), .q(v676obus), .dec(dec[676]));
wire [data_w*6-1:0] v677ibus;
wire [temp_w*6-1:0] v677obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU677 (.l(l[677*data_w +:data_w]), .r(v677ibus), .q(v677obus), .dec(dec[677]));
wire [data_w*6-1:0] v678ibus;
wire [temp_w*6-1:0] v678obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU678 (.l(l[678*data_w +:data_w]), .r(v678ibus), .q(v678obus), .dec(dec[678]));
wire [data_w*6-1:0] v679ibus;
wire [temp_w*6-1:0] v679obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU679 (.l(l[679*data_w +:data_w]), .r(v679ibus), .q(v679obus), .dec(dec[679]));
wire [data_w*6-1:0] v680ibus;
wire [temp_w*6-1:0] v680obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU680 (.l(l[680*data_w +:data_w]), .r(v680ibus), .q(v680obus), .dec(dec[680]));
wire [data_w*6-1:0] v681ibus;
wire [temp_w*6-1:0] v681obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU681 (.l(l[681*data_w +:data_w]), .r(v681ibus), .q(v681obus), .dec(dec[681]));
wire [data_w*6-1:0] v682ibus;
wire [temp_w*6-1:0] v682obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU682 (.l(l[682*data_w +:data_w]), .r(v682ibus), .q(v682obus), .dec(dec[682]));
wire [data_w*6-1:0] v683ibus;
wire [temp_w*6-1:0] v683obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU683 (.l(l[683*data_w +:data_w]), .r(v683ibus), .q(v683obus), .dec(dec[683]));
wire [data_w*6-1:0] v684ibus;
wire [temp_w*6-1:0] v684obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU684 (.l(l[684*data_w +:data_w]), .r(v684ibus), .q(v684obus), .dec(dec[684]));
wire [data_w*6-1:0] v685ibus;
wire [temp_w*6-1:0] v685obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU685 (.l(l[685*data_w +:data_w]), .r(v685ibus), .q(v685obus), .dec(dec[685]));
wire [data_w*6-1:0] v686ibus;
wire [temp_w*6-1:0] v686obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU686 (.l(l[686*data_w +:data_w]), .r(v686ibus), .q(v686obus), .dec(dec[686]));
wire [data_w*6-1:0] v687ibus;
wire [temp_w*6-1:0] v687obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU687 (.l(l[687*data_w +:data_w]), .r(v687ibus), .q(v687obus), .dec(dec[687]));
wire [data_w*6-1:0] v688ibus;
wire [temp_w*6-1:0] v688obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU688 (.l(l[688*data_w +:data_w]), .r(v688ibus), .q(v688obus), .dec(dec[688]));
wire [data_w*6-1:0] v689ibus;
wire [temp_w*6-1:0] v689obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU689 (.l(l[689*data_w +:data_w]), .r(v689ibus), .q(v689obus), .dec(dec[689]));
wire [data_w*6-1:0] v690ibus;
wire [temp_w*6-1:0] v690obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU690 (.l(l[690*data_w +:data_w]), .r(v690ibus), .q(v690obus), .dec(dec[690]));
wire [data_w*6-1:0] v691ibus;
wire [temp_w*6-1:0] v691obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU691 (.l(l[691*data_w +:data_w]), .r(v691ibus), .q(v691obus), .dec(dec[691]));
wire [data_w*6-1:0] v692ibus;
wire [temp_w*6-1:0] v692obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU692 (.l(l[692*data_w +:data_w]), .r(v692ibus), .q(v692obus), .dec(dec[692]));
wire [data_w*6-1:0] v693ibus;
wire [temp_w*6-1:0] v693obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU693 (.l(l[693*data_w +:data_w]), .r(v693ibus), .q(v693obus), .dec(dec[693]));
wire [data_w*6-1:0] v694ibus;
wire [temp_w*6-1:0] v694obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU694 (.l(l[694*data_w +:data_w]), .r(v694ibus), .q(v694obus), .dec(dec[694]));
wire [data_w*6-1:0] v695ibus;
wire [temp_w*6-1:0] v695obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU695 (.l(l[695*data_w +:data_w]), .r(v695ibus), .q(v695obus), .dec(dec[695]));
wire [data_w*6-1:0] v696ibus;
wire [temp_w*6-1:0] v696obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU696 (.l(l[696*data_w +:data_w]), .r(v696ibus), .q(v696obus), .dec(dec[696]));
wire [data_w*6-1:0] v697ibus;
wire [temp_w*6-1:0] v697obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU697 (.l(l[697*data_w +:data_w]), .r(v697ibus), .q(v697obus), .dec(dec[697]));
wire [data_w*6-1:0] v698ibus;
wire [temp_w*6-1:0] v698obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU698 (.l(l[698*data_w +:data_w]), .r(v698ibus), .q(v698obus), .dec(dec[698]));
wire [data_w*6-1:0] v699ibus;
wire [temp_w*6-1:0] v699obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU699 (.l(l[699*data_w +:data_w]), .r(v699ibus), .q(v699obus), .dec(dec[699]));
wire [data_w*6-1:0] v700ibus;
wire [temp_w*6-1:0] v700obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU700 (.l(l[700*data_w +:data_w]), .r(v700ibus), .q(v700obus), .dec(dec[700]));
wire [data_w*6-1:0] v701ibus;
wire [temp_w*6-1:0] v701obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU701 (.l(l[701*data_w +:data_w]), .r(v701ibus), .q(v701obus), .dec(dec[701]));
wire [data_w*6-1:0] v702ibus;
wire [temp_w*6-1:0] v702obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU702 (.l(l[702*data_w +:data_w]), .r(v702ibus), .q(v702obus), .dec(dec[702]));
wire [data_w*6-1:0] v703ibus;
wire [temp_w*6-1:0] v703obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU703 (.l(l[703*data_w +:data_w]), .r(v703ibus), .q(v703obus), .dec(dec[703]));
wire [data_w*6-1:0] v704ibus;
wire [temp_w*6-1:0] v704obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU704 (.l(l[704*data_w +:data_w]), .r(v704ibus), .q(v704obus), .dec(dec[704]));
wire [data_w*6-1:0] v705ibus;
wire [temp_w*6-1:0] v705obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU705 (.l(l[705*data_w +:data_w]), .r(v705ibus), .q(v705obus), .dec(dec[705]));
wire [data_w*6-1:0] v706ibus;
wire [temp_w*6-1:0] v706obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU706 (.l(l[706*data_w +:data_w]), .r(v706ibus), .q(v706obus), .dec(dec[706]));
wire [data_w*6-1:0] v707ibus;
wire [temp_w*6-1:0] v707obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU707 (.l(l[707*data_w +:data_w]), .r(v707ibus), .q(v707obus), .dec(dec[707]));
wire [data_w*6-1:0] v708ibus;
wire [temp_w*6-1:0] v708obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU708 (.l(l[708*data_w +:data_w]), .r(v708ibus), .q(v708obus), .dec(dec[708]));
wire [data_w*6-1:0] v709ibus;
wire [temp_w*6-1:0] v709obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU709 (.l(l[709*data_w +:data_w]), .r(v709ibus), .q(v709obus), .dec(dec[709]));
wire [data_w*6-1:0] v710ibus;
wire [temp_w*6-1:0] v710obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU710 (.l(l[710*data_w +:data_w]), .r(v710ibus), .q(v710obus), .dec(dec[710]));
wire [data_w*6-1:0] v711ibus;
wire [temp_w*6-1:0] v711obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU711 (.l(l[711*data_w +:data_w]), .r(v711ibus), .q(v711obus), .dec(dec[711]));
wire [data_w*6-1:0] v712ibus;
wire [temp_w*6-1:0] v712obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU712 (.l(l[712*data_w +:data_w]), .r(v712ibus), .q(v712obus), .dec(dec[712]));
wire [data_w*6-1:0] v713ibus;
wire [temp_w*6-1:0] v713obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU713 (.l(l[713*data_w +:data_w]), .r(v713ibus), .q(v713obus), .dec(dec[713]));
wire [data_w*6-1:0] v714ibus;
wire [temp_w*6-1:0] v714obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU714 (.l(l[714*data_w +:data_w]), .r(v714ibus), .q(v714obus), .dec(dec[714]));
wire [data_w*6-1:0] v715ibus;
wire [temp_w*6-1:0] v715obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU715 (.l(l[715*data_w +:data_w]), .r(v715ibus), .q(v715obus), .dec(dec[715]));
wire [data_w*6-1:0] v716ibus;
wire [temp_w*6-1:0] v716obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU716 (.l(l[716*data_w +:data_w]), .r(v716ibus), .q(v716obus), .dec(dec[716]));
wire [data_w*6-1:0] v717ibus;
wire [temp_w*6-1:0] v717obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU717 (.l(l[717*data_w +:data_w]), .r(v717ibus), .q(v717obus), .dec(dec[717]));
wire [data_w*6-1:0] v718ibus;
wire [temp_w*6-1:0] v718obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU718 (.l(l[718*data_w +:data_w]), .r(v718ibus), .q(v718obus), .dec(dec[718]));
wire [data_w*6-1:0] v719ibus;
wire [temp_w*6-1:0] v719obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU719 (.l(l[719*data_w +:data_w]), .r(v719ibus), .q(v719obus), .dec(dec[719]));
wire [data_w*6-1:0] v720ibus;
wire [temp_w*6-1:0] v720obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU720 (.l(l[720*data_w +:data_w]), .r(v720ibus), .q(v720obus), .dec(dec[720]));
wire [data_w*6-1:0] v721ibus;
wire [temp_w*6-1:0] v721obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU721 (.l(l[721*data_w +:data_w]), .r(v721ibus), .q(v721obus), .dec(dec[721]));
wire [data_w*6-1:0] v722ibus;
wire [temp_w*6-1:0] v722obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU722 (.l(l[722*data_w +:data_w]), .r(v722ibus), .q(v722obus), .dec(dec[722]));
wire [data_w*6-1:0] v723ibus;
wire [temp_w*6-1:0] v723obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU723 (.l(l[723*data_w +:data_w]), .r(v723ibus), .q(v723obus), .dec(dec[723]));
wire [data_w*6-1:0] v724ibus;
wire [temp_w*6-1:0] v724obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU724 (.l(l[724*data_w +:data_w]), .r(v724ibus), .q(v724obus), .dec(dec[724]));
wire [data_w*6-1:0] v725ibus;
wire [temp_w*6-1:0] v725obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU725 (.l(l[725*data_w +:data_w]), .r(v725ibus), .q(v725obus), .dec(dec[725]));
wire [data_w*6-1:0] v726ibus;
wire [temp_w*6-1:0] v726obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU726 (.l(l[726*data_w +:data_w]), .r(v726ibus), .q(v726obus), .dec(dec[726]));
wire [data_w*6-1:0] v727ibus;
wire [temp_w*6-1:0] v727obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU727 (.l(l[727*data_w +:data_w]), .r(v727ibus), .q(v727obus), .dec(dec[727]));
wire [data_w*6-1:0] v728ibus;
wire [temp_w*6-1:0] v728obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU728 (.l(l[728*data_w +:data_w]), .r(v728ibus), .q(v728obus), .dec(dec[728]));
wire [data_w*6-1:0] v729ibus;
wire [temp_w*6-1:0] v729obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU729 (.l(l[729*data_w +:data_w]), .r(v729ibus), .q(v729obus), .dec(dec[729]));
wire [data_w*6-1:0] v730ibus;
wire [temp_w*6-1:0] v730obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU730 (.l(l[730*data_w +:data_w]), .r(v730ibus), .q(v730obus), .dec(dec[730]));
wire [data_w*6-1:0] v731ibus;
wire [temp_w*6-1:0] v731obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU731 (.l(l[731*data_w +:data_w]), .r(v731ibus), .q(v731obus), .dec(dec[731]));
wire [data_w*6-1:0] v732ibus;
wire [temp_w*6-1:0] v732obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU732 (.l(l[732*data_w +:data_w]), .r(v732ibus), .q(v732obus), .dec(dec[732]));
wire [data_w*6-1:0] v733ibus;
wire [temp_w*6-1:0] v733obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU733 (.l(l[733*data_w +:data_w]), .r(v733ibus), .q(v733obus), .dec(dec[733]));
wire [data_w*6-1:0] v734ibus;
wire [temp_w*6-1:0] v734obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU734 (.l(l[734*data_w +:data_w]), .r(v734ibus), .q(v734obus), .dec(dec[734]));
wire [data_w*6-1:0] v735ibus;
wire [temp_w*6-1:0] v735obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU735 (.l(l[735*data_w +:data_w]), .r(v735ibus), .q(v735obus), .dec(dec[735]));
wire [data_w*6-1:0] v736ibus;
wire [temp_w*6-1:0] v736obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU736 (.l(l[736*data_w +:data_w]), .r(v736ibus), .q(v736obus), .dec(dec[736]));
wire [data_w*6-1:0] v737ibus;
wire [temp_w*6-1:0] v737obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU737 (.l(l[737*data_w +:data_w]), .r(v737ibus), .q(v737obus), .dec(dec[737]));
wire [data_w*6-1:0] v738ibus;
wire [temp_w*6-1:0] v738obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU738 (.l(l[738*data_w +:data_w]), .r(v738ibus), .q(v738obus), .dec(dec[738]));
wire [data_w*6-1:0] v739ibus;
wire [temp_w*6-1:0] v739obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU739 (.l(l[739*data_w +:data_w]), .r(v739ibus), .q(v739obus), .dec(dec[739]));
wire [data_w*6-1:0] v740ibus;
wire [temp_w*6-1:0] v740obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU740 (.l(l[740*data_w +:data_w]), .r(v740ibus), .q(v740obus), .dec(dec[740]));
wire [data_w*6-1:0] v741ibus;
wire [temp_w*6-1:0] v741obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU741 (.l(l[741*data_w +:data_w]), .r(v741ibus), .q(v741obus), .dec(dec[741]));
wire [data_w*6-1:0] v742ibus;
wire [temp_w*6-1:0] v742obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU742 (.l(l[742*data_w +:data_w]), .r(v742ibus), .q(v742obus), .dec(dec[742]));
wire [data_w*6-1:0] v743ibus;
wire [temp_w*6-1:0] v743obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU743 (.l(l[743*data_w +:data_w]), .r(v743ibus), .q(v743obus), .dec(dec[743]));
wire [data_w*6-1:0] v744ibus;
wire [temp_w*6-1:0] v744obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU744 (.l(l[744*data_w +:data_w]), .r(v744ibus), .q(v744obus), .dec(dec[744]));
wire [data_w*6-1:0] v745ibus;
wire [temp_w*6-1:0] v745obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU745 (.l(l[745*data_w +:data_w]), .r(v745ibus), .q(v745obus), .dec(dec[745]));
wire [data_w*6-1:0] v746ibus;
wire [temp_w*6-1:0] v746obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU746 (.l(l[746*data_w +:data_w]), .r(v746ibus), .q(v746obus), .dec(dec[746]));
wire [data_w*6-1:0] v747ibus;
wire [temp_w*6-1:0] v747obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU747 (.l(l[747*data_w +:data_w]), .r(v747ibus), .q(v747obus), .dec(dec[747]));
wire [data_w*6-1:0] v748ibus;
wire [temp_w*6-1:0] v748obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU748 (.l(l[748*data_w +:data_w]), .r(v748ibus), .q(v748obus), .dec(dec[748]));
wire [data_w*6-1:0] v749ibus;
wire [temp_w*6-1:0] v749obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU749 (.l(l[749*data_w +:data_w]), .r(v749ibus), .q(v749obus), .dec(dec[749]));
wire [data_w*6-1:0] v750ibus;
wire [temp_w*6-1:0] v750obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU750 (.l(l[750*data_w +:data_w]), .r(v750ibus), .q(v750obus), .dec(dec[750]));
wire [data_w*6-1:0] v751ibus;
wire [temp_w*6-1:0] v751obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU751 (.l(l[751*data_w +:data_w]), .r(v751ibus), .q(v751obus), .dec(dec[751]));
wire [data_w*6-1:0] v752ibus;
wire [temp_w*6-1:0] v752obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU752 (.l(l[752*data_w +:data_w]), .r(v752ibus), .q(v752obus), .dec(dec[752]));
wire [data_w*6-1:0] v753ibus;
wire [temp_w*6-1:0] v753obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU753 (.l(l[753*data_w +:data_w]), .r(v753ibus), .q(v753obus), .dec(dec[753]));
wire [data_w*6-1:0] v754ibus;
wire [temp_w*6-1:0] v754obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU754 (.l(l[754*data_w +:data_w]), .r(v754ibus), .q(v754obus), .dec(dec[754]));
wire [data_w*6-1:0] v755ibus;
wire [temp_w*6-1:0] v755obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU755 (.l(l[755*data_w +:data_w]), .r(v755ibus), .q(v755obus), .dec(dec[755]));
wire [data_w*6-1:0] v756ibus;
wire [temp_w*6-1:0] v756obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU756 (.l(l[756*data_w +:data_w]), .r(v756ibus), .q(v756obus), .dec(dec[756]));
wire [data_w*6-1:0] v757ibus;
wire [temp_w*6-1:0] v757obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU757 (.l(l[757*data_w +:data_w]), .r(v757ibus), .q(v757obus), .dec(dec[757]));
wire [data_w*6-1:0] v758ibus;
wire [temp_w*6-1:0] v758obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU758 (.l(l[758*data_w +:data_w]), .r(v758ibus), .q(v758obus), .dec(dec[758]));
wire [data_w*6-1:0] v759ibus;
wire [temp_w*6-1:0] v759obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU759 (.l(l[759*data_w +:data_w]), .r(v759ibus), .q(v759obus), .dec(dec[759]));
wire [data_w*6-1:0] v760ibus;
wire [temp_w*6-1:0] v760obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU760 (.l(l[760*data_w +:data_w]), .r(v760ibus), .q(v760obus), .dec(dec[760]));
wire [data_w*6-1:0] v761ibus;
wire [temp_w*6-1:0] v761obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU761 (.l(l[761*data_w +:data_w]), .r(v761ibus), .q(v761obus), .dec(dec[761]));
wire [data_w*6-1:0] v762ibus;
wire [temp_w*6-1:0] v762obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU762 (.l(l[762*data_w +:data_w]), .r(v762ibus), .q(v762obus), .dec(dec[762]));
wire [data_w*6-1:0] v763ibus;
wire [temp_w*6-1:0] v763obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU763 (.l(l[763*data_w +:data_w]), .r(v763ibus), .q(v763obus), .dec(dec[763]));
wire [data_w*6-1:0] v764ibus;
wire [temp_w*6-1:0] v764obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU764 (.l(l[764*data_w +:data_w]), .r(v764ibus), .q(v764obus), .dec(dec[764]));
wire [data_w*6-1:0] v765ibus;
wire [temp_w*6-1:0] v765obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU765 (.l(l[765*data_w +:data_w]), .r(v765ibus), .q(v765obus), .dec(dec[765]));
wire [data_w*6-1:0] v766ibus;
wire [temp_w*6-1:0] v766obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU766 (.l(l[766*data_w +:data_w]), .r(v766ibus), .q(v766obus), .dec(dec[766]));
wire [data_w*6-1:0] v767ibus;
wire [temp_w*6-1:0] v767obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU767 (.l(l[767*data_w +:data_w]), .r(v767ibus), .q(v767obus), .dec(dec[767]));
wire [data_w*3-1:0] v768ibus;
wire [temp_w*3-1:0] v768obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU768 (.l(l[768*data_w +:data_w]), .r(v768ibus), .q(v768obus), .dec(dec[768]));
wire [data_w*3-1:0] v769ibus;
wire [temp_w*3-1:0] v769obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU769 (.l(l[769*data_w +:data_w]), .r(v769ibus), .q(v769obus), .dec(dec[769]));
wire [data_w*3-1:0] v770ibus;
wire [temp_w*3-1:0] v770obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU770 (.l(l[770*data_w +:data_w]), .r(v770ibus), .q(v770obus), .dec(dec[770]));
wire [data_w*3-1:0] v771ibus;
wire [temp_w*3-1:0] v771obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU771 (.l(l[771*data_w +:data_w]), .r(v771ibus), .q(v771obus), .dec(dec[771]));
wire [data_w*3-1:0] v772ibus;
wire [temp_w*3-1:0] v772obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU772 (.l(l[772*data_w +:data_w]), .r(v772ibus), .q(v772obus), .dec(dec[772]));
wire [data_w*3-1:0] v773ibus;
wire [temp_w*3-1:0] v773obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU773 (.l(l[773*data_w +:data_w]), .r(v773ibus), .q(v773obus), .dec(dec[773]));
wire [data_w*3-1:0] v774ibus;
wire [temp_w*3-1:0] v774obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU774 (.l(l[774*data_w +:data_w]), .r(v774ibus), .q(v774obus), .dec(dec[774]));
wire [data_w*3-1:0] v775ibus;
wire [temp_w*3-1:0] v775obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU775 (.l(l[775*data_w +:data_w]), .r(v775ibus), .q(v775obus), .dec(dec[775]));
wire [data_w*3-1:0] v776ibus;
wire [temp_w*3-1:0] v776obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU776 (.l(l[776*data_w +:data_w]), .r(v776ibus), .q(v776obus), .dec(dec[776]));
wire [data_w*3-1:0] v777ibus;
wire [temp_w*3-1:0] v777obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU777 (.l(l[777*data_w +:data_w]), .r(v777ibus), .q(v777obus), .dec(dec[777]));
wire [data_w*3-1:0] v778ibus;
wire [temp_w*3-1:0] v778obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU778 (.l(l[778*data_w +:data_w]), .r(v778ibus), .q(v778obus), .dec(dec[778]));
wire [data_w*3-1:0] v779ibus;
wire [temp_w*3-1:0] v779obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU779 (.l(l[779*data_w +:data_w]), .r(v779ibus), .q(v779obus), .dec(dec[779]));
wire [data_w*3-1:0] v780ibus;
wire [temp_w*3-1:0] v780obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU780 (.l(l[780*data_w +:data_w]), .r(v780ibus), .q(v780obus), .dec(dec[780]));
wire [data_w*3-1:0] v781ibus;
wire [temp_w*3-1:0] v781obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU781 (.l(l[781*data_w +:data_w]), .r(v781ibus), .q(v781obus), .dec(dec[781]));
wire [data_w*3-1:0] v782ibus;
wire [temp_w*3-1:0] v782obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU782 (.l(l[782*data_w +:data_w]), .r(v782ibus), .q(v782obus), .dec(dec[782]));
wire [data_w*3-1:0] v783ibus;
wire [temp_w*3-1:0] v783obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU783 (.l(l[783*data_w +:data_w]), .r(v783ibus), .q(v783obus), .dec(dec[783]));
wire [data_w*3-1:0] v784ibus;
wire [temp_w*3-1:0] v784obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU784 (.l(l[784*data_w +:data_w]), .r(v784ibus), .q(v784obus), .dec(dec[784]));
wire [data_w*3-1:0] v785ibus;
wire [temp_w*3-1:0] v785obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU785 (.l(l[785*data_w +:data_w]), .r(v785ibus), .q(v785obus), .dec(dec[785]));
wire [data_w*3-1:0] v786ibus;
wire [temp_w*3-1:0] v786obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU786 (.l(l[786*data_w +:data_w]), .r(v786ibus), .q(v786obus), .dec(dec[786]));
wire [data_w*3-1:0] v787ibus;
wire [temp_w*3-1:0] v787obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU787 (.l(l[787*data_w +:data_w]), .r(v787ibus), .q(v787obus), .dec(dec[787]));
wire [data_w*3-1:0] v788ibus;
wire [temp_w*3-1:0] v788obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU788 (.l(l[788*data_w +:data_w]), .r(v788ibus), .q(v788obus), .dec(dec[788]));
wire [data_w*3-1:0] v789ibus;
wire [temp_w*3-1:0] v789obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU789 (.l(l[789*data_w +:data_w]), .r(v789ibus), .q(v789obus), .dec(dec[789]));
wire [data_w*3-1:0] v790ibus;
wire [temp_w*3-1:0] v790obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU790 (.l(l[790*data_w +:data_w]), .r(v790ibus), .q(v790obus), .dec(dec[790]));
wire [data_w*3-1:0] v791ibus;
wire [temp_w*3-1:0] v791obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU791 (.l(l[791*data_w +:data_w]), .r(v791ibus), .q(v791obus), .dec(dec[791]));
wire [data_w*3-1:0] v792ibus;
wire [temp_w*3-1:0] v792obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU792 (.l(l[792*data_w +:data_w]), .r(v792ibus), .q(v792obus), .dec(dec[792]));
wire [data_w*3-1:0] v793ibus;
wire [temp_w*3-1:0] v793obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU793 (.l(l[793*data_w +:data_w]), .r(v793ibus), .q(v793obus), .dec(dec[793]));
wire [data_w*3-1:0] v794ibus;
wire [temp_w*3-1:0] v794obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU794 (.l(l[794*data_w +:data_w]), .r(v794ibus), .q(v794obus), .dec(dec[794]));
wire [data_w*3-1:0] v795ibus;
wire [temp_w*3-1:0] v795obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU795 (.l(l[795*data_w +:data_w]), .r(v795ibus), .q(v795obus), .dec(dec[795]));
wire [data_w*3-1:0] v796ibus;
wire [temp_w*3-1:0] v796obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU796 (.l(l[796*data_w +:data_w]), .r(v796ibus), .q(v796obus), .dec(dec[796]));
wire [data_w*3-1:0] v797ibus;
wire [temp_w*3-1:0] v797obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU797 (.l(l[797*data_w +:data_w]), .r(v797ibus), .q(v797obus), .dec(dec[797]));
wire [data_w*3-1:0] v798ibus;
wire [temp_w*3-1:0] v798obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU798 (.l(l[798*data_w +:data_w]), .r(v798ibus), .q(v798obus), .dec(dec[798]));
wire [data_w*3-1:0] v799ibus;
wire [temp_w*3-1:0] v799obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU799 (.l(l[799*data_w +:data_w]), .r(v799ibus), .q(v799obus), .dec(dec[799]));
wire [data_w*3-1:0] v800ibus;
wire [temp_w*3-1:0] v800obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU800 (.l(l[800*data_w +:data_w]), .r(v800ibus), .q(v800obus), .dec(dec[800]));
wire [data_w*3-1:0] v801ibus;
wire [temp_w*3-1:0] v801obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU801 (.l(l[801*data_w +:data_w]), .r(v801ibus), .q(v801obus), .dec(dec[801]));
wire [data_w*3-1:0] v802ibus;
wire [temp_w*3-1:0] v802obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU802 (.l(l[802*data_w +:data_w]), .r(v802ibus), .q(v802obus), .dec(dec[802]));
wire [data_w*3-1:0] v803ibus;
wire [temp_w*3-1:0] v803obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU803 (.l(l[803*data_w +:data_w]), .r(v803ibus), .q(v803obus), .dec(dec[803]));
wire [data_w*3-1:0] v804ibus;
wire [temp_w*3-1:0] v804obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU804 (.l(l[804*data_w +:data_w]), .r(v804ibus), .q(v804obus), .dec(dec[804]));
wire [data_w*3-1:0] v805ibus;
wire [temp_w*3-1:0] v805obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU805 (.l(l[805*data_w +:data_w]), .r(v805ibus), .q(v805obus), .dec(dec[805]));
wire [data_w*3-1:0] v806ibus;
wire [temp_w*3-1:0] v806obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU806 (.l(l[806*data_w +:data_w]), .r(v806ibus), .q(v806obus), .dec(dec[806]));
wire [data_w*3-1:0] v807ibus;
wire [temp_w*3-1:0] v807obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU807 (.l(l[807*data_w +:data_w]), .r(v807ibus), .q(v807obus), .dec(dec[807]));
wire [data_w*3-1:0] v808ibus;
wire [temp_w*3-1:0] v808obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU808 (.l(l[808*data_w +:data_w]), .r(v808ibus), .q(v808obus), .dec(dec[808]));
wire [data_w*3-1:0] v809ibus;
wire [temp_w*3-1:0] v809obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU809 (.l(l[809*data_w +:data_w]), .r(v809ibus), .q(v809obus), .dec(dec[809]));
wire [data_w*3-1:0] v810ibus;
wire [temp_w*3-1:0] v810obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU810 (.l(l[810*data_w +:data_w]), .r(v810ibus), .q(v810obus), .dec(dec[810]));
wire [data_w*3-1:0] v811ibus;
wire [temp_w*3-1:0] v811obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU811 (.l(l[811*data_w +:data_w]), .r(v811ibus), .q(v811obus), .dec(dec[811]));
wire [data_w*3-1:0] v812ibus;
wire [temp_w*3-1:0] v812obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU812 (.l(l[812*data_w +:data_w]), .r(v812ibus), .q(v812obus), .dec(dec[812]));
wire [data_w*3-1:0] v813ibus;
wire [temp_w*3-1:0] v813obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU813 (.l(l[813*data_w +:data_w]), .r(v813ibus), .q(v813obus), .dec(dec[813]));
wire [data_w*3-1:0] v814ibus;
wire [temp_w*3-1:0] v814obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU814 (.l(l[814*data_w +:data_w]), .r(v814ibus), .q(v814obus), .dec(dec[814]));
wire [data_w*3-1:0] v815ibus;
wire [temp_w*3-1:0] v815obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU815 (.l(l[815*data_w +:data_w]), .r(v815ibus), .q(v815obus), .dec(dec[815]));
wire [data_w*3-1:0] v816ibus;
wire [temp_w*3-1:0] v816obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU816 (.l(l[816*data_w +:data_w]), .r(v816ibus), .q(v816obus), .dec(dec[816]));
wire [data_w*3-1:0] v817ibus;
wire [temp_w*3-1:0] v817obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU817 (.l(l[817*data_w +:data_w]), .r(v817ibus), .q(v817obus), .dec(dec[817]));
wire [data_w*3-1:0] v818ibus;
wire [temp_w*3-1:0] v818obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU818 (.l(l[818*data_w +:data_w]), .r(v818ibus), .q(v818obus), .dec(dec[818]));
wire [data_w*3-1:0] v819ibus;
wire [temp_w*3-1:0] v819obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU819 (.l(l[819*data_w +:data_w]), .r(v819ibus), .q(v819obus), .dec(dec[819]));
wire [data_w*3-1:0] v820ibus;
wire [temp_w*3-1:0] v820obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU820 (.l(l[820*data_w +:data_w]), .r(v820ibus), .q(v820obus), .dec(dec[820]));
wire [data_w*3-1:0] v821ibus;
wire [temp_w*3-1:0] v821obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU821 (.l(l[821*data_w +:data_w]), .r(v821ibus), .q(v821obus), .dec(dec[821]));
wire [data_w*3-1:0] v822ibus;
wire [temp_w*3-1:0] v822obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU822 (.l(l[822*data_w +:data_w]), .r(v822ibus), .q(v822obus), .dec(dec[822]));
wire [data_w*3-1:0] v823ibus;
wire [temp_w*3-1:0] v823obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU823 (.l(l[823*data_w +:data_w]), .r(v823ibus), .q(v823obus), .dec(dec[823]));
wire [data_w*3-1:0] v824ibus;
wire [temp_w*3-1:0] v824obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU824 (.l(l[824*data_w +:data_w]), .r(v824ibus), .q(v824obus), .dec(dec[824]));
wire [data_w*3-1:0] v825ibus;
wire [temp_w*3-1:0] v825obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU825 (.l(l[825*data_w +:data_w]), .r(v825ibus), .q(v825obus), .dec(dec[825]));
wire [data_w*3-1:0] v826ibus;
wire [temp_w*3-1:0] v826obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU826 (.l(l[826*data_w +:data_w]), .r(v826ibus), .q(v826obus), .dec(dec[826]));
wire [data_w*3-1:0] v827ibus;
wire [temp_w*3-1:0] v827obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU827 (.l(l[827*data_w +:data_w]), .r(v827ibus), .q(v827obus), .dec(dec[827]));
wire [data_w*3-1:0] v828ibus;
wire [temp_w*3-1:0] v828obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU828 (.l(l[828*data_w +:data_w]), .r(v828ibus), .q(v828obus), .dec(dec[828]));
wire [data_w*3-1:0] v829ibus;
wire [temp_w*3-1:0] v829obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU829 (.l(l[829*data_w +:data_w]), .r(v829ibus), .q(v829obus), .dec(dec[829]));
wire [data_w*3-1:0] v830ibus;
wire [temp_w*3-1:0] v830obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU830 (.l(l[830*data_w +:data_w]), .r(v830ibus), .q(v830obus), .dec(dec[830]));
wire [data_w*3-1:0] v831ibus;
wire [temp_w*3-1:0] v831obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU831 (.l(l[831*data_w +:data_w]), .r(v831ibus), .q(v831obus), .dec(dec[831]));
wire [data_w*3-1:0] v832ibus;
wire [temp_w*3-1:0] v832obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU832 (.l(l[832*data_w +:data_w]), .r(v832ibus), .q(v832obus), .dec(dec[832]));
wire [data_w*3-1:0] v833ibus;
wire [temp_w*3-1:0] v833obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU833 (.l(l[833*data_w +:data_w]), .r(v833ibus), .q(v833obus), .dec(dec[833]));
wire [data_w*3-1:0] v834ibus;
wire [temp_w*3-1:0] v834obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU834 (.l(l[834*data_w +:data_w]), .r(v834ibus), .q(v834obus), .dec(dec[834]));
wire [data_w*3-1:0] v835ibus;
wire [temp_w*3-1:0] v835obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU835 (.l(l[835*data_w +:data_w]), .r(v835ibus), .q(v835obus), .dec(dec[835]));
wire [data_w*3-1:0] v836ibus;
wire [temp_w*3-1:0] v836obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU836 (.l(l[836*data_w +:data_w]), .r(v836ibus), .q(v836obus), .dec(dec[836]));
wire [data_w*3-1:0] v837ibus;
wire [temp_w*3-1:0] v837obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU837 (.l(l[837*data_w +:data_w]), .r(v837ibus), .q(v837obus), .dec(dec[837]));
wire [data_w*3-1:0] v838ibus;
wire [temp_w*3-1:0] v838obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU838 (.l(l[838*data_w +:data_w]), .r(v838ibus), .q(v838obus), .dec(dec[838]));
wire [data_w*3-1:0] v839ibus;
wire [temp_w*3-1:0] v839obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU839 (.l(l[839*data_w +:data_w]), .r(v839ibus), .q(v839obus), .dec(dec[839]));
wire [data_w*3-1:0] v840ibus;
wire [temp_w*3-1:0] v840obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU840 (.l(l[840*data_w +:data_w]), .r(v840ibus), .q(v840obus), .dec(dec[840]));
wire [data_w*3-1:0] v841ibus;
wire [temp_w*3-1:0] v841obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU841 (.l(l[841*data_w +:data_w]), .r(v841ibus), .q(v841obus), .dec(dec[841]));
wire [data_w*3-1:0] v842ibus;
wire [temp_w*3-1:0] v842obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU842 (.l(l[842*data_w +:data_w]), .r(v842ibus), .q(v842obus), .dec(dec[842]));
wire [data_w*3-1:0] v843ibus;
wire [temp_w*3-1:0] v843obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU843 (.l(l[843*data_w +:data_w]), .r(v843ibus), .q(v843obus), .dec(dec[843]));
wire [data_w*3-1:0] v844ibus;
wire [temp_w*3-1:0] v844obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU844 (.l(l[844*data_w +:data_w]), .r(v844ibus), .q(v844obus), .dec(dec[844]));
wire [data_w*3-1:0] v845ibus;
wire [temp_w*3-1:0] v845obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU845 (.l(l[845*data_w +:data_w]), .r(v845ibus), .q(v845obus), .dec(dec[845]));
wire [data_w*3-1:0] v846ibus;
wire [temp_w*3-1:0] v846obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU846 (.l(l[846*data_w +:data_w]), .r(v846ibus), .q(v846obus), .dec(dec[846]));
wire [data_w*3-1:0] v847ibus;
wire [temp_w*3-1:0] v847obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU847 (.l(l[847*data_w +:data_w]), .r(v847ibus), .q(v847obus), .dec(dec[847]));
wire [data_w*3-1:0] v848ibus;
wire [temp_w*3-1:0] v848obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU848 (.l(l[848*data_w +:data_w]), .r(v848ibus), .q(v848obus), .dec(dec[848]));
wire [data_w*3-1:0] v849ibus;
wire [temp_w*3-1:0] v849obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU849 (.l(l[849*data_w +:data_w]), .r(v849ibus), .q(v849obus), .dec(dec[849]));
wire [data_w*3-1:0] v850ibus;
wire [temp_w*3-1:0] v850obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU850 (.l(l[850*data_w +:data_w]), .r(v850ibus), .q(v850obus), .dec(dec[850]));
wire [data_w*3-1:0] v851ibus;
wire [temp_w*3-1:0] v851obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU851 (.l(l[851*data_w +:data_w]), .r(v851ibus), .q(v851obus), .dec(dec[851]));
wire [data_w*3-1:0] v852ibus;
wire [temp_w*3-1:0] v852obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU852 (.l(l[852*data_w +:data_w]), .r(v852ibus), .q(v852obus), .dec(dec[852]));
wire [data_w*3-1:0] v853ibus;
wire [temp_w*3-1:0] v853obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU853 (.l(l[853*data_w +:data_w]), .r(v853ibus), .q(v853obus), .dec(dec[853]));
wire [data_w*3-1:0] v854ibus;
wire [temp_w*3-1:0] v854obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU854 (.l(l[854*data_w +:data_w]), .r(v854ibus), .q(v854obus), .dec(dec[854]));
wire [data_w*3-1:0] v855ibus;
wire [temp_w*3-1:0] v855obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU855 (.l(l[855*data_w +:data_w]), .r(v855ibus), .q(v855obus), .dec(dec[855]));
wire [data_w*3-1:0] v856ibus;
wire [temp_w*3-1:0] v856obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU856 (.l(l[856*data_w +:data_w]), .r(v856ibus), .q(v856obus), .dec(dec[856]));
wire [data_w*3-1:0] v857ibus;
wire [temp_w*3-1:0] v857obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU857 (.l(l[857*data_w +:data_w]), .r(v857ibus), .q(v857obus), .dec(dec[857]));
wire [data_w*3-1:0] v858ibus;
wire [temp_w*3-1:0] v858obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU858 (.l(l[858*data_w +:data_w]), .r(v858ibus), .q(v858obus), .dec(dec[858]));
wire [data_w*3-1:0] v859ibus;
wire [temp_w*3-1:0] v859obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU859 (.l(l[859*data_w +:data_w]), .r(v859ibus), .q(v859obus), .dec(dec[859]));
wire [data_w*3-1:0] v860ibus;
wire [temp_w*3-1:0] v860obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU860 (.l(l[860*data_w +:data_w]), .r(v860ibus), .q(v860obus), .dec(dec[860]));
wire [data_w*3-1:0] v861ibus;
wire [temp_w*3-1:0] v861obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU861 (.l(l[861*data_w +:data_w]), .r(v861ibus), .q(v861obus), .dec(dec[861]));
wire [data_w*3-1:0] v862ibus;
wire [temp_w*3-1:0] v862obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU862 (.l(l[862*data_w +:data_w]), .r(v862ibus), .q(v862obus), .dec(dec[862]));
wire [data_w*3-1:0] v863ibus;
wire [temp_w*3-1:0] v863obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU863 (.l(l[863*data_w +:data_w]), .r(v863ibus), .q(v863obus), .dec(dec[863]));
wire [data_w*6-1:0] v864ibus;
wire [temp_w*6-1:0] v864obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU864 (.l(l[864*data_w +:data_w]), .r(v864ibus), .q(v864obus), .dec(dec[864]));
wire [data_w*6-1:0] v865ibus;
wire [temp_w*6-1:0] v865obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU865 (.l(l[865*data_w +:data_w]), .r(v865ibus), .q(v865obus), .dec(dec[865]));
wire [data_w*6-1:0] v866ibus;
wire [temp_w*6-1:0] v866obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU866 (.l(l[866*data_w +:data_w]), .r(v866ibus), .q(v866obus), .dec(dec[866]));
wire [data_w*6-1:0] v867ibus;
wire [temp_w*6-1:0] v867obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU867 (.l(l[867*data_w +:data_w]), .r(v867ibus), .q(v867obus), .dec(dec[867]));
wire [data_w*6-1:0] v868ibus;
wire [temp_w*6-1:0] v868obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU868 (.l(l[868*data_w +:data_w]), .r(v868ibus), .q(v868obus), .dec(dec[868]));
wire [data_w*6-1:0] v869ibus;
wire [temp_w*6-1:0] v869obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU869 (.l(l[869*data_w +:data_w]), .r(v869ibus), .q(v869obus), .dec(dec[869]));
wire [data_w*6-1:0] v870ibus;
wire [temp_w*6-1:0] v870obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU870 (.l(l[870*data_w +:data_w]), .r(v870ibus), .q(v870obus), .dec(dec[870]));
wire [data_w*6-1:0] v871ibus;
wire [temp_w*6-1:0] v871obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU871 (.l(l[871*data_w +:data_w]), .r(v871ibus), .q(v871obus), .dec(dec[871]));
wire [data_w*6-1:0] v872ibus;
wire [temp_w*6-1:0] v872obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU872 (.l(l[872*data_w +:data_w]), .r(v872ibus), .q(v872obus), .dec(dec[872]));
wire [data_w*6-1:0] v873ibus;
wire [temp_w*6-1:0] v873obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU873 (.l(l[873*data_w +:data_w]), .r(v873ibus), .q(v873obus), .dec(dec[873]));
wire [data_w*6-1:0] v874ibus;
wire [temp_w*6-1:0] v874obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU874 (.l(l[874*data_w +:data_w]), .r(v874ibus), .q(v874obus), .dec(dec[874]));
wire [data_w*6-1:0] v875ibus;
wire [temp_w*6-1:0] v875obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU875 (.l(l[875*data_w +:data_w]), .r(v875ibus), .q(v875obus), .dec(dec[875]));
wire [data_w*6-1:0] v876ibus;
wire [temp_w*6-1:0] v876obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU876 (.l(l[876*data_w +:data_w]), .r(v876ibus), .q(v876obus), .dec(dec[876]));
wire [data_w*6-1:0] v877ibus;
wire [temp_w*6-1:0] v877obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU877 (.l(l[877*data_w +:data_w]), .r(v877ibus), .q(v877obus), .dec(dec[877]));
wire [data_w*6-1:0] v878ibus;
wire [temp_w*6-1:0] v878obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU878 (.l(l[878*data_w +:data_w]), .r(v878ibus), .q(v878obus), .dec(dec[878]));
wire [data_w*6-1:0] v879ibus;
wire [temp_w*6-1:0] v879obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU879 (.l(l[879*data_w +:data_w]), .r(v879ibus), .q(v879obus), .dec(dec[879]));
wire [data_w*6-1:0] v880ibus;
wire [temp_w*6-1:0] v880obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU880 (.l(l[880*data_w +:data_w]), .r(v880ibus), .q(v880obus), .dec(dec[880]));
wire [data_w*6-1:0] v881ibus;
wire [temp_w*6-1:0] v881obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU881 (.l(l[881*data_w +:data_w]), .r(v881ibus), .q(v881obus), .dec(dec[881]));
wire [data_w*6-1:0] v882ibus;
wire [temp_w*6-1:0] v882obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU882 (.l(l[882*data_w +:data_w]), .r(v882ibus), .q(v882obus), .dec(dec[882]));
wire [data_w*6-1:0] v883ibus;
wire [temp_w*6-1:0] v883obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU883 (.l(l[883*data_w +:data_w]), .r(v883ibus), .q(v883obus), .dec(dec[883]));
wire [data_w*6-1:0] v884ibus;
wire [temp_w*6-1:0] v884obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU884 (.l(l[884*data_w +:data_w]), .r(v884ibus), .q(v884obus), .dec(dec[884]));
wire [data_w*6-1:0] v885ibus;
wire [temp_w*6-1:0] v885obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU885 (.l(l[885*data_w +:data_w]), .r(v885ibus), .q(v885obus), .dec(dec[885]));
wire [data_w*6-1:0] v886ibus;
wire [temp_w*6-1:0] v886obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU886 (.l(l[886*data_w +:data_w]), .r(v886ibus), .q(v886obus), .dec(dec[886]));
wire [data_w*6-1:0] v887ibus;
wire [temp_w*6-1:0] v887obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU887 (.l(l[887*data_w +:data_w]), .r(v887ibus), .q(v887obus), .dec(dec[887]));
wire [data_w*6-1:0] v888ibus;
wire [temp_w*6-1:0] v888obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU888 (.l(l[888*data_w +:data_w]), .r(v888ibus), .q(v888obus), .dec(dec[888]));
wire [data_w*6-1:0] v889ibus;
wire [temp_w*6-1:0] v889obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU889 (.l(l[889*data_w +:data_w]), .r(v889ibus), .q(v889obus), .dec(dec[889]));
wire [data_w*6-1:0] v890ibus;
wire [temp_w*6-1:0] v890obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU890 (.l(l[890*data_w +:data_w]), .r(v890ibus), .q(v890obus), .dec(dec[890]));
wire [data_w*6-1:0] v891ibus;
wire [temp_w*6-1:0] v891obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU891 (.l(l[891*data_w +:data_w]), .r(v891ibus), .q(v891obus), .dec(dec[891]));
wire [data_w*6-1:0] v892ibus;
wire [temp_w*6-1:0] v892obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU892 (.l(l[892*data_w +:data_w]), .r(v892ibus), .q(v892obus), .dec(dec[892]));
wire [data_w*6-1:0] v893ibus;
wire [temp_w*6-1:0] v893obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU893 (.l(l[893*data_w +:data_w]), .r(v893ibus), .q(v893obus), .dec(dec[893]));
wire [data_w*6-1:0] v894ibus;
wire [temp_w*6-1:0] v894obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU894 (.l(l[894*data_w +:data_w]), .r(v894ibus), .q(v894obus), .dec(dec[894]));
wire [data_w*6-1:0] v895ibus;
wire [temp_w*6-1:0] v895obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU895 (.l(l[895*data_w +:data_w]), .r(v895ibus), .q(v895obus), .dec(dec[895]));
wire [data_w*6-1:0] v896ibus;
wire [temp_w*6-1:0] v896obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU896 (.l(l[896*data_w +:data_w]), .r(v896ibus), .q(v896obus), .dec(dec[896]));
wire [data_w*6-1:0] v897ibus;
wire [temp_w*6-1:0] v897obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU897 (.l(l[897*data_w +:data_w]), .r(v897ibus), .q(v897obus), .dec(dec[897]));
wire [data_w*6-1:0] v898ibus;
wire [temp_w*6-1:0] v898obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU898 (.l(l[898*data_w +:data_w]), .r(v898ibus), .q(v898obus), .dec(dec[898]));
wire [data_w*6-1:0] v899ibus;
wire [temp_w*6-1:0] v899obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU899 (.l(l[899*data_w +:data_w]), .r(v899ibus), .q(v899obus), .dec(dec[899]));
wire [data_w*6-1:0] v900ibus;
wire [temp_w*6-1:0] v900obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU900 (.l(l[900*data_w +:data_w]), .r(v900ibus), .q(v900obus), .dec(dec[900]));
wire [data_w*6-1:0] v901ibus;
wire [temp_w*6-1:0] v901obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU901 (.l(l[901*data_w +:data_w]), .r(v901ibus), .q(v901obus), .dec(dec[901]));
wire [data_w*6-1:0] v902ibus;
wire [temp_w*6-1:0] v902obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU902 (.l(l[902*data_w +:data_w]), .r(v902ibus), .q(v902obus), .dec(dec[902]));
wire [data_w*6-1:0] v903ibus;
wire [temp_w*6-1:0] v903obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU903 (.l(l[903*data_w +:data_w]), .r(v903ibus), .q(v903obus), .dec(dec[903]));
wire [data_w*6-1:0] v904ibus;
wire [temp_w*6-1:0] v904obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU904 (.l(l[904*data_w +:data_w]), .r(v904ibus), .q(v904obus), .dec(dec[904]));
wire [data_w*6-1:0] v905ibus;
wire [temp_w*6-1:0] v905obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU905 (.l(l[905*data_w +:data_w]), .r(v905ibus), .q(v905obus), .dec(dec[905]));
wire [data_w*6-1:0] v906ibus;
wire [temp_w*6-1:0] v906obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU906 (.l(l[906*data_w +:data_w]), .r(v906ibus), .q(v906obus), .dec(dec[906]));
wire [data_w*6-1:0] v907ibus;
wire [temp_w*6-1:0] v907obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU907 (.l(l[907*data_w +:data_w]), .r(v907ibus), .q(v907obus), .dec(dec[907]));
wire [data_w*6-1:0] v908ibus;
wire [temp_w*6-1:0] v908obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU908 (.l(l[908*data_w +:data_w]), .r(v908ibus), .q(v908obus), .dec(dec[908]));
wire [data_w*6-1:0] v909ibus;
wire [temp_w*6-1:0] v909obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU909 (.l(l[909*data_w +:data_w]), .r(v909ibus), .q(v909obus), .dec(dec[909]));
wire [data_w*6-1:0] v910ibus;
wire [temp_w*6-1:0] v910obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU910 (.l(l[910*data_w +:data_w]), .r(v910ibus), .q(v910obus), .dec(dec[910]));
wire [data_w*6-1:0] v911ibus;
wire [temp_w*6-1:0] v911obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU911 (.l(l[911*data_w +:data_w]), .r(v911ibus), .q(v911obus), .dec(dec[911]));
wire [data_w*6-1:0] v912ibus;
wire [temp_w*6-1:0] v912obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU912 (.l(l[912*data_w +:data_w]), .r(v912ibus), .q(v912obus), .dec(dec[912]));
wire [data_w*6-1:0] v913ibus;
wire [temp_w*6-1:0] v913obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU913 (.l(l[913*data_w +:data_w]), .r(v913ibus), .q(v913obus), .dec(dec[913]));
wire [data_w*6-1:0] v914ibus;
wire [temp_w*6-1:0] v914obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU914 (.l(l[914*data_w +:data_w]), .r(v914ibus), .q(v914obus), .dec(dec[914]));
wire [data_w*6-1:0] v915ibus;
wire [temp_w*6-1:0] v915obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU915 (.l(l[915*data_w +:data_w]), .r(v915ibus), .q(v915obus), .dec(dec[915]));
wire [data_w*6-1:0] v916ibus;
wire [temp_w*6-1:0] v916obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU916 (.l(l[916*data_w +:data_w]), .r(v916ibus), .q(v916obus), .dec(dec[916]));
wire [data_w*6-1:0] v917ibus;
wire [temp_w*6-1:0] v917obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU917 (.l(l[917*data_w +:data_w]), .r(v917ibus), .q(v917obus), .dec(dec[917]));
wire [data_w*6-1:0] v918ibus;
wire [temp_w*6-1:0] v918obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU918 (.l(l[918*data_w +:data_w]), .r(v918ibus), .q(v918obus), .dec(dec[918]));
wire [data_w*6-1:0] v919ibus;
wire [temp_w*6-1:0] v919obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU919 (.l(l[919*data_w +:data_w]), .r(v919ibus), .q(v919obus), .dec(dec[919]));
wire [data_w*6-1:0] v920ibus;
wire [temp_w*6-1:0] v920obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU920 (.l(l[920*data_w +:data_w]), .r(v920ibus), .q(v920obus), .dec(dec[920]));
wire [data_w*6-1:0] v921ibus;
wire [temp_w*6-1:0] v921obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU921 (.l(l[921*data_w +:data_w]), .r(v921ibus), .q(v921obus), .dec(dec[921]));
wire [data_w*6-1:0] v922ibus;
wire [temp_w*6-1:0] v922obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU922 (.l(l[922*data_w +:data_w]), .r(v922ibus), .q(v922obus), .dec(dec[922]));
wire [data_w*6-1:0] v923ibus;
wire [temp_w*6-1:0] v923obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU923 (.l(l[923*data_w +:data_w]), .r(v923ibus), .q(v923obus), .dec(dec[923]));
wire [data_w*6-1:0] v924ibus;
wire [temp_w*6-1:0] v924obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU924 (.l(l[924*data_w +:data_w]), .r(v924ibus), .q(v924obus), .dec(dec[924]));
wire [data_w*6-1:0] v925ibus;
wire [temp_w*6-1:0] v925obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU925 (.l(l[925*data_w +:data_w]), .r(v925ibus), .q(v925obus), .dec(dec[925]));
wire [data_w*6-1:0] v926ibus;
wire [temp_w*6-1:0] v926obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU926 (.l(l[926*data_w +:data_w]), .r(v926ibus), .q(v926obus), .dec(dec[926]));
wire [data_w*6-1:0] v927ibus;
wire [temp_w*6-1:0] v927obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU927 (.l(l[927*data_w +:data_w]), .r(v927ibus), .q(v927obus), .dec(dec[927]));
wire [data_w*6-1:0] v928ibus;
wire [temp_w*6-1:0] v928obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU928 (.l(l[928*data_w +:data_w]), .r(v928ibus), .q(v928obus), .dec(dec[928]));
wire [data_w*6-1:0] v929ibus;
wire [temp_w*6-1:0] v929obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU929 (.l(l[929*data_w +:data_w]), .r(v929ibus), .q(v929obus), .dec(dec[929]));
wire [data_w*6-1:0] v930ibus;
wire [temp_w*6-1:0] v930obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU930 (.l(l[930*data_w +:data_w]), .r(v930ibus), .q(v930obus), .dec(dec[930]));
wire [data_w*6-1:0] v931ibus;
wire [temp_w*6-1:0] v931obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU931 (.l(l[931*data_w +:data_w]), .r(v931ibus), .q(v931obus), .dec(dec[931]));
wire [data_w*6-1:0] v932ibus;
wire [temp_w*6-1:0] v932obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU932 (.l(l[932*data_w +:data_w]), .r(v932ibus), .q(v932obus), .dec(dec[932]));
wire [data_w*6-1:0] v933ibus;
wire [temp_w*6-1:0] v933obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU933 (.l(l[933*data_w +:data_w]), .r(v933ibus), .q(v933obus), .dec(dec[933]));
wire [data_w*6-1:0] v934ibus;
wire [temp_w*6-1:0] v934obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU934 (.l(l[934*data_w +:data_w]), .r(v934ibus), .q(v934obus), .dec(dec[934]));
wire [data_w*6-1:0] v935ibus;
wire [temp_w*6-1:0] v935obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU935 (.l(l[935*data_w +:data_w]), .r(v935ibus), .q(v935obus), .dec(dec[935]));
wire [data_w*6-1:0] v936ibus;
wire [temp_w*6-1:0] v936obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU936 (.l(l[936*data_w +:data_w]), .r(v936ibus), .q(v936obus), .dec(dec[936]));
wire [data_w*6-1:0] v937ibus;
wire [temp_w*6-1:0] v937obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU937 (.l(l[937*data_w +:data_w]), .r(v937ibus), .q(v937obus), .dec(dec[937]));
wire [data_w*6-1:0] v938ibus;
wire [temp_w*6-1:0] v938obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU938 (.l(l[938*data_w +:data_w]), .r(v938ibus), .q(v938obus), .dec(dec[938]));
wire [data_w*6-1:0] v939ibus;
wire [temp_w*6-1:0] v939obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU939 (.l(l[939*data_w +:data_w]), .r(v939ibus), .q(v939obus), .dec(dec[939]));
wire [data_w*6-1:0] v940ibus;
wire [temp_w*6-1:0] v940obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU940 (.l(l[940*data_w +:data_w]), .r(v940ibus), .q(v940obus), .dec(dec[940]));
wire [data_w*6-1:0] v941ibus;
wire [temp_w*6-1:0] v941obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU941 (.l(l[941*data_w +:data_w]), .r(v941ibus), .q(v941obus), .dec(dec[941]));
wire [data_w*6-1:0] v942ibus;
wire [temp_w*6-1:0] v942obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU942 (.l(l[942*data_w +:data_w]), .r(v942ibus), .q(v942obus), .dec(dec[942]));
wire [data_w*6-1:0] v943ibus;
wire [temp_w*6-1:0] v943obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU943 (.l(l[943*data_w +:data_w]), .r(v943ibus), .q(v943obus), .dec(dec[943]));
wire [data_w*6-1:0] v944ibus;
wire [temp_w*6-1:0] v944obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU944 (.l(l[944*data_w +:data_w]), .r(v944ibus), .q(v944obus), .dec(dec[944]));
wire [data_w*6-1:0] v945ibus;
wire [temp_w*6-1:0] v945obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU945 (.l(l[945*data_w +:data_w]), .r(v945ibus), .q(v945obus), .dec(dec[945]));
wire [data_w*6-1:0] v946ibus;
wire [temp_w*6-1:0] v946obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU946 (.l(l[946*data_w +:data_w]), .r(v946ibus), .q(v946obus), .dec(dec[946]));
wire [data_w*6-1:0] v947ibus;
wire [temp_w*6-1:0] v947obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU947 (.l(l[947*data_w +:data_w]), .r(v947ibus), .q(v947obus), .dec(dec[947]));
wire [data_w*6-1:0] v948ibus;
wire [temp_w*6-1:0] v948obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU948 (.l(l[948*data_w +:data_w]), .r(v948ibus), .q(v948obus), .dec(dec[948]));
wire [data_w*6-1:0] v949ibus;
wire [temp_w*6-1:0] v949obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU949 (.l(l[949*data_w +:data_w]), .r(v949ibus), .q(v949obus), .dec(dec[949]));
wire [data_w*6-1:0] v950ibus;
wire [temp_w*6-1:0] v950obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU950 (.l(l[950*data_w +:data_w]), .r(v950ibus), .q(v950obus), .dec(dec[950]));
wire [data_w*6-1:0] v951ibus;
wire [temp_w*6-1:0] v951obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU951 (.l(l[951*data_w +:data_w]), .r(v951ibus), .q(v951obus), .dec(dec[951]));
wire [data_w*6-1:0] v952ibus;
wire [temp_w*6-1:0] v952obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU952 (.l(l[952*data_w +:data_w]), .r(v952ibus), .q(v952obus), .dec(dec[952]));
wire [data_w*6-1:0] v953ibus;
wire [temp_w*6-1:0] v953obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU953 (.l(l[953*data_w +:data_w]), .r(v953ibus), .q(v953obus), .dec(dec[953]));
wire [data_w*6-1:0] v954ibus;
wire [temp_w*6-1:0] v954obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU954 (.l(l[954*data_w +:data_w]), .r(v954ibus), .q(v954obus), .dec(dec[954]));
wire [data_w*6-1:0] v955ibus;
wire [temp_w*6-1:0] v955obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU955 (.l(l[955*data_w +:data_w]), .r(v955ibus), .q(v955obus), .dec(dec[955]));
wire [data_w*6-1:0] v956ibus;
wire [temp_w*6-1:0] v956obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU956 (.l(l[956*data_w +:data_w]), .r(v956ibus), .q(v956obus), .dec(dec[956]));
wire [data_w*6-1:0] v957ibus;
wire [temp_w*6-1:0] v957obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU957 (.l(l[957*data_w +:data_w]), .r(v957ibus), .q(v957obus), .dec(dec[957]));
wire [data_w*6-1:0] v958ibus;
wire [temp_w*6-1:0] v958obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU958 (.l(l[958*data_w +:data_w]), .r(v958ibus), .q(v958obus), .dec(dec[958]));
wire [data_w*6-1:0] v959ibus;
wire [temp_w*6-1:0] v959obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU959 (.l(l[959*data_w +:data_w]), .r(v959ibus), .q(v959obus), .dec(dec[959]));
wire [data_w*3-1:0] v960ibus;
wire [temp_w*3-1:0] v960obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU960 (.l(l[960*data_w +:data_w]), .r(v960ibus), .q(v960obus), .dec(dec[960]));
wire [data_w*3-1:0] v961ibus;
wire [temp_w*3-1:0] v961obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU961 (.l(l[961*data_w +:data_w]), .r(v961ibus), .q(v961obus), .dec(dec[961]));
wire [data_w*3-1:0] v962ibus;
wire [temp_w*3-1:0] v962obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU962 (.l(l[962*data_w +:data_w]), .r(v962ibus), .q(v962obus), .dec(dec[962]));
wire [data_w*3-1:0] v963ibus;
wire [temp_w*3-1:0] v963obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU963 (.l(l[963*data_w +:data_w]), .r(v963ibus), .q(v963obus), .dec(dec[963]));
wire [data_w*3-1:0] v964ibus;
wire [temp_w*3-1:0] v964obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU964 (.l(l[964*data_w +:data_w]), .r(v964ibus), .q(v964obus), .dec(dec[964]));
wire [data_w*3-1:0] v965ibus;
wire [temp_w*3-1:0] v965obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU965 (.l(l[965*data_w +:data_w]), .r(v965ibus), .q(v965obus), .dec(dec[965]));
wire [data_w*3-1:0] v966ibus;
wire [temp_w*3-1:0] v966obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU966 (.l(l[966*data_w +:data_w]), .r(v966ibus), .q(v966obus), .dec(dec[966]));
wire [data_w*3-1:0] v967ibus;
wire [temp_w*3-1:0] v967obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU967 (.l(l[967*data_w +:data_w]), .r(v967ibus), .q(v967obus), .dec(dec[967]));
wire [data_w*3-1:0] v968ibus;
wire [temp_w*3-1:0] v968obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU968 (.l(l[968*data_w +:data_w]), .r(v968ibus), .q(v968obus), .dec(dec[968]));
wire [data_w*3-1:0] v969ibus;
wire [temp_w*3-1:0] v969obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU969 (.l(l[969*data_w +:data_w]), .r(v969ibus), .q(v969obus), .dec(dec[969]));
wire [data_w*3-1:0] v970ibus;
wire [temp_w*3-1:0] v970obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU970 (.l(l[970*data_w +:data_w]), .r(v970ibus), .q(v970obus), .dec(dec[970]));
wire [data_w*3-1:0] v971ibus;
wire [temp_w*3-1:0] v971obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU971 (.l(l[971*data_w +:data_w]), .r(v971ibus), .q(v971obus), .dec(dec[971]));
wire [data_w*3-1:0] v972ibus;
wire [temp_w*3-1:0] v972obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU972 (.l(l[972*data_w +:data_w]), .r(v972ibus), .q(v972obus), .dec(dec[972]));
wire [data_w*3-1:0] v973ibus;
wire [temp_w*3-1:0] v973obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU973 (.l(l[973*data_w +:data_w]), .r(v973ibus), .q(v973obus), .dec(dec[973]));
wire [data_w*3-1:0] v974ibus;
wire [temp_w*3-1:0] v974obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU974 (.l(l[974*data_w +:data_w]), .r(v974ibus), .q(v974obus), .dec(dec[974]));
wire [data_w*3-1:0] v975ibus;
wire [temp_w*3-1:0] v975obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU975 (.l(l[975*data_w +:data_w]), .r(v975ibus), .q(v975obus), .dec(dec[975]));
wire [data_w*3-1:0] v976ibus;
wire [temp_w*3-1:0] v976obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU976 (.l(l[976*data_w +:data_w]), .r(v976ibus), .q(v976obus), .dec(dec[976]));
wire [data_w*3-1:0] v977ibus;
wire [temp_w*3-1:0] v977obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU977 (.l(l[977*data_w +:data_w]), .r(v977ibus), .q(v977obus), .dec(dec[977]));
wire [data_w*3-1:0] v978ibus;
wire [temp_w*3-1:0] v978obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU978 (.l(l[978*data_w +:data_w]), .r(v978ibus), .q(v978obus), .dec(dec[978]));
wire [data_w*3-1:0] v979ibus;
wire [temp_w*3-1:0] v979obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU979 (.l(l[979*data_w +:data_w]), .r(v979ibus), .q(v979obus), .dec(dec[979]));
wire [data_w*3-1:0] v980ibus;
wire [temp_w*3-1:0] v980obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU980 (.l(l[980*data_w +:data_w]), .r(v980ibus), .q(v980obus), .dec(dec[980]));
wire [data_w*3-1:0] v981ibus;
wire [temp_w*3-1:0] v981obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU981 (.l(l[981*data_w +:data_w]), .r(v981ibus), .q(v981obus), .dec(dec[981]));
wire [data_w*3-1:0] v982ibus;
wire [temp_w*3-1:0] v982obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU982 (.l(l[982*data_w +:data_w]), .r(v982ibus), .q(v982obus), .dec(dec[982]));
wire [data_w*3-1:0] v983ibus;
wire [temp_w*3-1:0] v983obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU983 (.l(l[983*data_w +:data_w]), .r(v983ibus), .q(v983obus), .dec(dec[983]));
wire [data_w*3-1:0] v984ibus;
wire [temp_w*3-1:0] v984obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU984 (.l(l[984*data_w +:data_w]), .r(v984ibus), .q(v984obus), .dec(dec[984]));
wire [data_w*3-1:0] v985ibus;
wire [temp_w*3-1:0] v985obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU985 (.l(l[985*data_w +:data_w]), .r(v985ibus), .q(v985obus), .dec(dec[985]));
wire [data_w*3-1:0] v986ibus;
wire [temp_w*3-1:0] v986obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU986 (.l(l[986*data_w +:data_w]), .r(v986ibus), .q(v986obus), .dec(dec[986]));
wire [data_w*3-1:0] v987ibus;
wire [temp_w*3-1:0] v987obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU987 (.l(l[987*data_w +:data_w]), .r(v987ibus), .q(v987obus), .dec(dec[987]));
wire [data_w*3-1:0] v988ibus;
wire [temp_w*3-1:0] v988obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU988 (.l(l[988*data_w +:data_w]), .r(v988ibus), .q(v988obus), .dec(dec[988]));
wire [data_w*3-1:0] v989ibus;
wire [temp_w*3-1:0] v989obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU989 (.l(l[989*data_w +:data_w]), .r(v989ibus), .q(v989obus), .dec(dec[989]));
wire [data_w*3-1:0] v990ibus;
wire [temp_w*3-1:0] v990obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU990 (.l(l[990*data_w +:data_w]), .r(v990ibus), .q(v990obus), .dec(dec[990]));
wire [data_w*3-1:0] v991ibus;
wire [temp_w*3-1:0] v991obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU991 (.l(l[991*data_w +:data_w]), .r(v991ibus), .q(v991obus), .dec(dec[991]));
wire [data_w*3-1:0] v992ibus;
wire [temp_w*3-1:0] v992obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU992 (.l(l[992*data_w +:data_w]), .r(v992ibus), .q(v992obus), .dec(dec[992]));
wire [data_w*3-1:0] v993ibus;
wire [temp_w*3-1:0] v993obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU993 (.l(l[993*data_w +:data_w]), .r(v993ibus), .q(v993obus), .dec(dec[993]));
wire [data_w*3-1:0] v994ibus;
wire [temp_w*3-1:0] v994obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU994 (.l(l[994*data_w +:data_w]), .r(v994ibus), .q(v994obus), .dec(dec[994]));
wire [data_w*3-1:0] v995ibus;
wire [temp_w*3-1:0] v995obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU995 (.l(l[995*data_w +:data_w]), .r(v995ibus), .q(v995obus), .dec(dec[995]));
wire [data_w*3-1:0] v996ibus;
wire [temp_w*3-1:0] v996obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU996 (.l(l[996*data_w +:data_w]), .r(v996ibus), .q(v996obus), .dec(dec[996]));
wire [data_w*3-1:0] v997ibus;
wire [temp_w*3-1:0] v997obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU997 (.l(l[997*data_w +:data_w]), .r(v997ibus), .q(v997obus), .dec(dec[997]));
wire [data_w*3-1:0] v998ibus;
wire [temp_w*3-1:0] v998obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU998 (.l(l[998*data_w +:data_w]), .r(v998ibus), .q(v998obus), .dec(dec[998]));
wire [data_w*3-1:0] v999ibus;
wire [temp_w*3-1:0] v999obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU999 (.l(l[999*data_w +:data_w]), .r(v999ibus), .q(v999obus), .dec(dec[999]));
wire [data_w*3-1:0] v1000ibus;
wire [temp_w*3-1:0] v1000obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1000 (.l(l[1000*data_w +:data_w]), .r(v1000ibus), .q(v1000obus), .dec(dec[1000]));
wire [data_w*3-1:0] v1001ibus;
wire [temp_w*3-1:0] v1001obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1001 (.l(l[1001*data_w +:data_w]), .r(v1001ibus), .q(v1001obus), .dec(dec[1001]));
wire [data_w*3-1:0] v1002ibus;
wire [temp_w*3-1:0] v1002obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1002 (.l(l[1002*data_w +:data_w]), .r(v1002ibus), .q(v1002obus), .dec(dec[1002]));
wire [data_w*3-1:0] v1003ibus;
wire [temp_w*3-1:0] v1003obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1003 (.l(l[1003*data_w +:data_w]), .r(v1003ibus), .q(v1003obus), .dec(dec[1003]));
wire [data_w*3-1:0] v1004ibus;
wire [temp_w*3-1:0] v1004obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1004 (.l(l[1004*data_w +:data_w]), .r(v1004ibus), .q(v1004obus), .dec(dec[1004]));
wire [data_w*3-1:0] v1005ibus;
wire [temp_w*3-1:0] v1005obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1005 (.l(l[1005*data_w +:data_w]), .r(v1005ibus), .q(v1005obus), .dec(dec[1005]));
wire [data_w*3-1:0] v1006ibus;
wire [temp_w*3-1:0] v1006obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1006 (.l(l[1006*data_w +:data_w]), .r(v1006ibus), .q(v1006obus), .dec(dec[1006]));
wire [data_w*3-1:0] v1007ibus;
wire [temp_w*3-1:0] v1007obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1007 (.l(l[1007*data_w +:data_w]), .r(v1007ibus), .q(v1007obus), .dec(dec[1007]));
wire [data_w*3-1:0] v1008ibus;
wire [temp_w*3-1:0] v1008obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1008 (.l(l[1008*data_w +:data_w]), .r(v1008ibus), .q(v1008obus), .dec(dec[1008]));
wire [data_w*3-1:0] v1009ibus;
wire [temp_w*3-1:0] v1009obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1009 (.l(l[1009*data_w +:data_w]), .r(v1009ibus), .q(v1009obus), .dec(dec[1009]));
wire [data_w*3-1:0] v1010ibus;
wire [temp_w*3-1:0] v1010obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1010 (.l(l[1010*data_w +:data_w]), .r(v1010ibus), .q(v1010obus), .dec(dec[1010]));
wire [data_w*3-1:0] v1011ibus;
wire [temp_w*3-1:0] v1011obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1011 (.l(l[1011*data_w +:data_w]), .r(v1011ibus), .q(v1011obus), .dec(dec[1011]));
wire [data_w*3-1:0] v1012ibus;
wire [temp_w*3-1:0] v1012obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1012 (.l(l[1012*data_w +:data_w]), .r(v1012ibus), .q(v1012obus), .dec(dec[1012]));
wire [data_w*3-1:0] v1013ibus;
wire [temp_w*3-1:0] v1013obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1013 (.l(l[1013*data_w +:data_w]), .r(v1013ibus), .q(v1013obus), .dec(dec[1013]));
wire [data_w*3-1:0] v1014ibus;
wire [temp_w*3-1:0] v1014obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1014 (.l(l[1014*data_w +:data_w]), .r(v1014ibus), .q(v1014obus), .dec(dec[1014]));
wire [data_w*3-1:0] v1015ibus;
wire [temp_w*3-1:0] v1015obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1015 (.l(l[1015*data_w +:data_w]), .r(v1015ibus), .q(v1015obus), .dec(dec[1015]));
wire [data_w*3-1:0] v1016ibus;
wire [temp_w*3-1:0] v1016obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1016 (.l(l[1016*data_w +:data_w]), .r(v1016ibus), .q(v1016obus), .dec(dec[1016]));
wire [data_w*3-1:0] v1017ibus;
wire [temp_w*3-1:0] v1017obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1017 (.l(l[1017*data_w +:data_w]), .r(v1017ibus), .q(v1017obus), .dec(dec[1017]));
wire [data_w*3-1:0] v1018ibus;
wire [temp_w*3-1:0] v1018obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1018 (.l(l[1018*data_w +:data_w]), .r(v1018ibus), .q(v1018obus), .dec(dec[1018]));
wire [data_w*3-1:0] v1019ibus;
wire [temp_w*3-1:0] v1019obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1019 (.l(l[1019*data_w +:data_w]), .r(v1019ibus), .q(v1019obus), .dec(dec[1019]));
wire [data_w*3-1:0] v1020ibus;
wire [temp_w*3-1:0] v1020obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1020 (.l(l[1020*data_w +:data_w]), .r(v1020ibus), .q(v1020obus), .dec(dec[1020]));
wire [data_w*3-1:0] v1021ibus;
wire [temp_w*3-1:0] v1021obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1021 (.l(l[1021*data_w +:data_w]), .r(v1021ibus), .q(v1021obus), .dec(dec[1021]));
wire [data_w*3-1:0] v1022ibus;
wire [temp_w*3-1:0] v1022obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1022 (.l(l[1022*data_w +:data_w]), .r(v1022ibus), .q(v1022obus), .dec(dec[1022]));
wire [data_w*3-1:0] v1023ibus;
wire [temp_w*3-1:0] v1023obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1023 (.l(l[1023*data_w +:data_w]), .r(v1023ibus), .q(v1023obus), .dec(dec[1023]));
wire [data_w*3-1:0] v1024ibus;
wire [temp_w*3-1:0] v1024obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1024 (.l(l[1024*data_w +:data_w]), .r(v1024ibus), .q(v1024obus), .dec(dec[1024]));
wire [data_w*3-1:0] v1025ibus;
wire [temp_w*3-1:0] v1025obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1025 (.l(l[1025*data_w +:data_w]), .r(v1025ibus), .q(v1025obus), .dec(dec[1025]));
wire [data_w*3-1:0] v1026ibus;
wire [temp_w*3-1:0] v1026obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1026 (.l(l[1026*data_w +:data_w]), .r(v1026ibus), .q(v1026obus), .dec(dec[1026]));
wire [data_w*3-1:0] v1027ibus;
wire [temp_w*3-1:0] v1027obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1027 (.l(l[1027*data_w +:data_w]), .r(v1027ibus), .q(v1027obus), .dec(dec[1027]));
wire [data_w*3-1:0] v1028ibus;
wire [temp_w*3-1:0] v1028obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1028 (.l(l[1028*data_w +:data_w]), .r(v1028ibus), .q(v1028obus), .dec(dec[1028]));
wire [data_w*3-1:0] v1029ibus;
wire [temp_w*3-1:0] v1029obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1029 (.l(l[1029*data_w +:data_w]), .r(v1029ibus), .q(v1029obus), .dec(dec[1029]));
wire [data_w*3-1:0] v1030ibus;
wire [temp_w*3-1:0] v1030obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1030 (.l(l[1030*data_w +:data_w]), .r(v1030ibus), .q(v1030obus), .dec(dec[1030]));
wire [data_w*3-1:0] v1031ibus;
wire [temp_w*3-1:0] v1031obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1031 (.l(l[1031*data_w +:data_w]), .r(v1031ibus), .q(v1031obus), .dec(dec[1031]));
wire [data_w*3-1:0] v1032ibus;
wire [temp_w*3-1:0] v1032obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1032 (.l(l[1032*data_w +:data_w]), .r(v1032ibus), .q(v1032obus), .dec(dec[1032]));
wire [data_w*3-1:0] v1033ibus;
wire [temp_w*3-1:0] v1033obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1033 (.l(l[1033*data_w +:data_w]), .r(v1033ibus), .q(v1033obus), .dec(dec[1033]));
wire [data_w*3-1:0] v1034ibus;
wire [temp_w*3-1:0] v1034obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1034 (.l(l[1034*data_w +:data_w]), .r(v1034ibus), .q(v1034obus), .dec(dec[1034]));
wire [data_w*3-1:0] v1035ibus;
wire [temp_w*3-1:0] v1035obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1035 (.l(l[1035*data_w +:data_w]), .r(v1035ibus), .q(v1035obus), .dec(dec[1035]));
wire [data_w*3-1:0] v1036ibus;
wire [temp_w*3-1:0] v1036obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1036 (.l(l[1036*data_w +:data_w]), .r(v1036ibus), .q(v1036obus), .dec(dec[1036]));
wire [data_w*3-1:0] v1037ibus;
wire [temp_w*3-1:0] v1037obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1037 (.l(l[1037*data_w +:data_w]), .r(v1037ibus), .q(v1037obus), .dec(dec[1037]));
wire [data_w*3-1:0] v1038ibus;
wire [temp_w*3-1:0] v1038obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1038 (.l(l[1038*data_w +:data_w]), .r(v1038ibus), .q(v1038obus), .dec(dec[1038]));
wire [data_w*3-1:0] v1039ibus;
wire [temp_w*3-1:0] v1039obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1039 (.l(l[1039*data_w +:data_w]), .r(v1039ibus), .q(v1039obus), .dec(dec[1039]));
wire [data_w*3-1:0] v1040ibus;
wire [temp_w*3-1:0] v1040obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1040 (.l(l[1040*data_w +:data_w]), .r(v1040ibus), .q(v1040obus), .dec(dec[1040]));
wire [data_w*3-1:0] v1041ibus;
wire [temp_w*3-1:0] v1041obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1041 (.l(l[1041*data_w +:data_w]), .r(v1041ibus), .q(v1041obus), .dec(dec[1041]));
wire [data_w*3-1:0] v1042ibus;
wire [temp_w*3-1:0] v1042obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1042 (.l(l[1042*data_w +:data_w]), .r(v1042ibus), .q(v1042obus), .dec(dec[1042]));
wire [data_w*3-1:0] v1043ibus;
wire [temp_w*3-1:0] v1043obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1043 (.l(l[1043*data_w +:data_w]), .r(v1043ibus), .q(v1043obus), .dec(dec[1043]));
wire [data_w*3-1:0] v1044ibus;
wire [temp_w*3-1:0] v1044obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1044 (.l(l[1044*data_w +:data_w]), .r(v1044ibus), .q(v1044obus), .dec(dec[1044]));
wire [data_w*3-1:0] v1045ibus;
wire [temp_w*3-1:0] v1045obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1045 (.l(l[1045*data_w +:data_w]), .r(v1045ibus), .q(v1045obus), .dec(dec[1045]));
wire [data_w*3-1:0] v1046ibus;
wire [temp_w*3-1:0] v1046obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1046 (.l(l[1046*data_w +:data_w]), .r(v1046ibus), .q(v1046obus), .dec(dec[1046]));
wire [data_w*3-1:0] v1047ibus;
wire [temp_w*3-1:0] v1047obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1047 (.l(l[1047*data_w +:data_w]), .r(v1047ibus), .q(v1047obus), .dec(dec[1047]));
wire [data_w*3-1:0] v1048ibus;
wire [temp_w*3-1:0] v1048obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1048 (.l(l[1048*data_w +:data_w]), .r(v1048ibus), .q(v1048obus), .dec(dec[1048]));
wire [data_w*3-1:0] v1049ibus;
wire [temp_w*3-1:0] v1049obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1049 (.l(l[1049*data_w +:data_w]), .r(v1049ibus), .q(v1049obus), .dec(dec[1049]));
wire [data_w*3-1:0] v1050ibus;
wire [temp_w*3-1:0] v1050obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1050 (.l(l[1050*data_w +:data_w]), .r(v1050ibus), .q(v1050obus), .dec(dec[1050]));
wire [data_w*3-1:0] v1051ibus;
wire [temp_w*3-1:0] v1051obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1051 (.l(l[1051*data_w +:data_w]), .r(v1051ibus), .q(v1051obus), .dec(dec[1051]));
wire [data_w*3-1:0] v1052ibus;
wire [temp_w*3-1:0] v1052obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1052 (.l(l[1052*data_w +:data_w]), .r(v1052ibus), .q(v1052obus), .dec(dec[1052]));
wire [data_w*3-1:0] v1053ibus;
wire [temp_w*3-1:0] v1053obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1053 (.l(l[1053*data_w +:data_w]), .r(v1053ibus), .q(v1053obus), .dec(dec[1053]));
wire [data_w*3-1:0] v1054ibus;
wire [temp_w*3-1:0] v1054obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1054 (.l(l[1054*data_w +:data_w]), .r(v1054ibus), .q(v1054obus), .dec(dec[1054]));
wire [data_w*3-1:0] v1055ibus;
wire [temp_w*3-1:0] v1055obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1055 (.l(l[1055*data_w +:data_w]), .r(v1055ibus), .q(v1055obus), .dec(dec[1055]));
wire [data_w*6-1:0] v1056ibus;
wire [temp_w*6-1:0] v1056obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1056 (.l(l[1056*data_w +:data_w]), .r(v1056ibus), .q(v1056obus), .dec(dec[1056]));
wire [data_w*6-1:0] v1057ibus;
wire [temp_w*6-1:0] v1057obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1057 (.l(l[1057*data_w +:data_w]), .r(v1057ibus), .q(v1057obus), .dec(dec[1057]));
wire [data_w*6-1:0] v1058ibus;
wire [temp_w*6-1:0] v1058obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1058 (.l(l[1058*data_w +:data_w]), .r(v1058ibus), .q(v1058obus), .dec(dec[1058]));
wire [data_w*6-1:0] v1059ibus;
wire [temp_w*6-1:0] v1059obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1059 (.l(l[1059*data_w +:data_w]), .r(v1059ibus), .q(v1059obus), .dec(dec[1059]));
wire [data_w*6-1:0] v1060ibus;
wire [temp_w*6-1:0] v1060obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1060 (.l(l[1060*data_w +:data_w]), .r(v1060ibus), .q(v1060obus), .dec(dec[1060]));
wire [data_w*6-1:0] v1061ibus;
wire [temp_w*6-1:0] v1061obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1061 (.l(l[1061*data_w +:data_w]), .r(v1061ibus), .q(v1061obus), .dec(dec[1061]));
wire [data_w*6-1:0] v1062ibus;
wire [temp_w*6-1:0] v1062obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1062 (.l(l[1062*data_w +:data_w]), .r(v1062ibus), .q(v1062obus), .dec(dec[1062]));
wire [data_w*6-1:0] v1063ibus;
wire [temp_w*6-1:0] v1063obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1063 (.l(l[1063*data_w +:data_w]), .r(v1063ibus), .q(v1063obus), .dec(dec[1063]));
wire [data_w*6-1:0] v1064ibus;
wire [temp_w*6-1:0] v1064obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1064 (.l(l[1064*data_w +:data_w]), .r(v1064ibus), .q(v1064obus), .dec(dec[1064]));
wire [data_w*6-1:0] v1065ibus;
wire [temp_w*6-1:0] v1065obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1065 (.l(l[1065*data_w +:data_w]), .r(v1065ibus), .q(v1065obus), .dec(dec[1065]));
wire [data_w*6-1:0] v1066ibus;
wire [temp_w*6-1:0] v1066obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1066 (.l(l[1066*data_w +:data_w]), .r(v1066ibus), .q(v1066obus), .dec(dec[1066]));
wire [data_w*6-1:0] v1067ibus;
wire [temp_w*6-1:0] v1067obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1067 (.l(l[1067*data_w +:data_w]), .r(v1067ibus), .q(v1067obus), .dec(dec[1067]));
wire [data_w*6-1:0] v1068ibus;
wire [temp_w*6-1:0] v1068obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1068 (.l(l[1068*data_w +:data_w]), .r(v1068ibus), .q(v1068obus), .dec(dec[1068]));
wire [data_w*6-1:0] v1069ibus;
wire [temp_w*6-1:0] v1069obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1069 (.l(l[1069*data_w +:data_w]), .r(v1069ibus), .q(v1069obus), .dec(dec[1069]));
wire [data_w*6-1:0] v1070ibus;
wire [temp_w*6-1:0] v1070obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1070 (.l(l[1070*data_w +:data_w]), .r(v1070ibus), .q(v1070obus), .dec(dec[1070]));
wire [data_w*6-1:0] v1071ibus;
wire [temp_w*6-1:0] v1071obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1071 (.l(l[1071*data_w +:data_w]), .r(v1071ibus), .q(v1071obus), .dec(dec[1071]));
wire [data_w*6-1:0] v1072ibus;
wire [temp_w*6-1:0] v1072obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1072 (.l(l[1072*data_w +:data_w]), .r(v1072ibus), .q(v1072obus), .dec(dec[1072]));
wire [data_w*6-1:0] v1073ibus;
wire [temp_w*6-1:0] v1073obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1073 (.l(l[1073*data_w +:data_w]), .r(v1073ibus), .q(v1073obus), .dec(dec[1073]));
wire [data_w*6-1:0] v1074ibus;
wire [temp_w*6-1:0] v1074obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1074 (.l(l[1074*data_w +:data_w]), .r(v1074ibus), .q(v1074obus), .dec(dec[1074]));
wire [data_w*6-1:0] v1075ibus;
wire [temp_w*6-1:0] v1075obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1075 (.l(l[1075*data_w +:data_w]), .r(v1075ibus), .q(v1075obus), .dec(dec[1075]));
wire [data_w*6-1:0] v1076ibus;
wire [temp_w*6-1:0] v1076obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1076 (.l(l[1076*data_w +:data_w]), .r(v1076ibus), .q(v1076obus), .dec(dec[1076]));
wire [data_w*6-1:0] v1077ibus;
wire [temp_w*6-1:0] v1077obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1077 (.l(l[1077*data_w +:data_w]), .r(v1077ibus), .q(v1077obus), .dec(dec[1077]));
wire [data_w*6-1:0] v1078ibus;
wire [temp_w*6-1:0] v1078obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1078 (.l(l[1078*data_w +:data_w]), .r(v1078ibus), .q(v1078obus), .dec(dec[1078]));
wire [data_w*6-1:0] v1079ibus;
wire [temp_w*6-1:0] v1079obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1079 (.l(l[1079*data_w +:data_w]), .r(v1079ibus), .q(v1079obus), .dec(dec[1079]));
wire [data_w*6-1:0] v1080ibus;
wire [temp_w*6-1:0] v1080obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1080 (.l(l[1080*data_w +:data_w]), .r(v1080ibus), .q(v1080obus), .dec(dec[1080]));
wire [data_w*6-1:0] v1081ibus;
wire [temp_w*6-1:0] v1081obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1081 (.l(l[1081*data_w +:data_w]), .r(v1081ibus), .q(v1081obus), .dec(dec[1081]));
wire [data_w*6-1:0] v1082ibus;
wire [temp_w*6-1:0] v1082obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1082 (.l(l[1082*data_w +:data_w]), .r(v1082ibus), .q(v1082obus), .dec(dec[1082]));
wire [data_w*6-1:0] v1083ibus;
wire [temp_w*6-1:0] v1083obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1083 (.l(l[1083*data_w +:data_w]), .r(v1083ibus), .q(v1083obus), .dec(dec[1083]));
wire [data_w*6-1:0] v1084ibus;
wire [temp_w*6-1:0] v1084obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1084 (.l(l[1084*data_w +:data_w]), .r(v1084ibus), .q(v1084obus), .dec(dec[1084]));
wire [data_w*6-1:0] v1085ibus;
wire [temp_w*6-1:0] v1085obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1085 (.l(l[1085*data_w +:data_w]), .r(v1085ibus), .q(v1085obus), .dec(dec[1085]));
wire [data_w*6-1:0] v1086ibus;
wire [temp_w*6-1:0] v1086obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1086 (.l(l[1086*data_w +:data_w]), .r(v1086ibus), .q(v1086obus), .dec(dec[1086]));
wire [data_w*6-1:0] v1087ibus;
wire [temp_w*6-1:0] v1087obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1087 (.l(l[1087*data_w +:data_w]), .r(v1087ibus), .q(v1087obus), .dec(dec[1087]));
wire [data_w*6-1:0] v1088ibus;
wire [temp_w*6-1:0] v1088obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1088 (.l(l[1088*data_w +:data_w]), .r(v1088ibus), .q(v1088obus), .dec(dec[1088]));
wire [data_w*6-1:0] v1089ibus;
wire [temp_w*6-1:0] v1089obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1089 (.l(l[1089*data_w +:data_w]), .r(v1089ibus), .q(v1089obus), .dec(dec[1089]));
wire [data_w*6-1:0] v1090ibus;
wire [temp_w*6-1:0] v1090obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1090 (.l(l[1090*data_w +:data_w]), .r(v1090ibus), .q(v1090obus), .dec(dec[1090]));
wire [data_w*6-1:0] v1091ibus;
wire [temp_w*6-1:0] v1091obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1091 (.l(l[1091*data_w +:data_w]), .r(v1091ibus), .q(v1091obus), .dec(dec[1091]));
wire [data_w*6-1:0] v1092ibus;
wire [temp_w*6-1:0] v1092obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1092 (.l(l[1092*data_w +:data_w]), .r(v1092ibus), .q(v1092obus), .dec(dec[1092]));
wire [data_w*6-1:0] v1093ibus;
wire [temp_w*6-1:0] v1093obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1093 (.l(l[1093*data_w +:data_w]), .r(v1093ibus), .q(v1093obus), .dec(dec[1093]));
wire [data_w*6-1:0] v1094ibus;
wire [temp_w*6-1:0] v1094obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1094 (.l(l[1094*data_w +:data_w]), .r(v1094ibus), .q(v1094obus), .dec(dec[1094]));
wire [data_w*6-1:0] v1095ibus;
wire [temp_w*6-1:0] v1095obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1095 (.l(l[1095*data_w +:data_w]), .r(v1095ibus), .q(v1095obus), .dec(dec[1095]));
wire [data_w*6-1:0] v1096ibus;
wire [temp_w*6-1:0] v1096obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1096 (.l(l[1096*data_w +:data_w]), .r(v1096ibus), .q(v1096obus), .dec(dec[1096]));
wire [data_w*6-1:0] v1097ibus;
wire [temp_w*6-1:0] v1097obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1097 (.l(l[1097*data_w +:data_w]), .r(v1097ibus), .q(v1097obus), .dec(dec[1097]));
wire [data_w*6-1:0] v1098ibus;
wire [temp_w*6-1:0] v1098obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1098 (.l(l[1098*data_w +:data_w]), .r(v1098ibus), .q(v1098obus), .dec(dec[1098]));
wire [data_w*6-1:0] v1099ibus;
wire [temp_w*6-1:0] v1099obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1099 (.l(l[1099*data_w +:data_w]), .r(v1099ibus), .q(v1099obus), .dec(dec[1099]));
wire [data_w*6-1:0] v1100ibus;
wire [temp_w*6-1:0] v1100obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1100 (.l(l[1100*data_w +:data_w]), .r(v1100ibus), .q(v1100obus), .dec(dec[1100]));
wire [data_w*6-1:0] v1101ibus;
wire [temp_w*6-1:0] v1101obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1101 (.l(l[1101*data_w +:data_w]), .r(v1101ibus), .q(v1101obus), .dec(dec[1101]));
wire [data_w*6-1:0] v1102ibus;
wire [temp_w*6-1:0] v1102obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1102 (.l(l[1102*data_w +:data_w]), .r(v1102ibus), .q(v1102obus), .dec(dec[1102]));
wire [data_w*6-1:0] v1103ibus;
wire [temp_w*6-1:0] v1103obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1103 (.l(l[1103*data_w +:data_w]), .r(v1103ibus), .q(v1103obus), .dec(dec[1103]));
wire [data_w*6-1:0] v1104ibus;
wire [temp_w*6-1:0] v1104obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1104 (.l(l[1104*data_w +:data_w]), .r(v1104ibus), .q(v1104obus), .dec(dec[1104]));
wire [data_w*6-1:0] v1105ibus;
wire [temp_w*6-1:0] v1105obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1105 (.l(l[1105*data_w +:data_w]), .r(v1105ibus), .q(v1105obus), .dec(dec[1105]));
wire [data_w*6-1:0] v1106ibus;
wire [temp_w*6-1:0] v1106obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1106 (.l(l[1106*data_w +:data_w]), .r(v1106ibus), .q(v1106obus), .dec(dec[1106]));
wire [data_w*6-1:0] v1107ibus;
wire [temp_w*6-1:0] v1107obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1107 (.l(l[1107*data_w +:data_w]), .r(v1107ibus), .q(v1107obus), .dec(dec[1107]));
wire [data_w*6-1:0] v1108ibus;
wire [temp_w*6-1:0] v1108obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1108 (.l(l[1108*data_w +:data_w]), .r(v1108ibus), .q(v1108obus), .dec(dec[1108]));
wire [data_w*6-1:0] v1109ibus;
wire [temp_w*6-1:0] v1109obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1109 (.l(l[1109*data_w +:data_w]), .r(v1109ibus), .q(v1109obus), .dec(dec[1109]));
wire [data_w*6-1:0] v1110ibus;
wire [temp_w*6-1:0] v1110obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1110 (.l(l[1110*data_w +:data_w]), .r(v1110ibus), .q(v1110obus), .dec(dec[1110]));
wire [data_w*6-1:0] v1111ibus;
wire [temp_w*6-1:0] v1111obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1111 (.l(l[1111*data_w +:data_w]), .r(v1111ibus), .q(v1111obus), .dec(dec[1111]));
wire [data_w*6-1:0] v1112ibus;
wire [temp_w*6-1:0] v1112obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1112 (.l(l[1112*data_w +:data_w]), .r(v1112ibus), .q(v1112obus), .dec(dec[1112]));
wire [data_w*6-1:0] v1113ibus;
wire [temp_w*6-1:0] v1113obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1113 (.l(l[1113*data_w +:data_w]), .r(v1113ibus), .q(v1113obus), .dec(dec[1113]));
wire [data_w*6-1:0] v1114ibus;
wire [temp_w*6-1:0] v1114obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1114 (.l(l[1114*data_w +:data_w]), .r(v1114ibus), .q(v1114obus), .dec(dec[1114]));
wire [data_w*6-1:0] v1115ibus;
wire [temp_w*6-1:0] v1115obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1115 (.l(l[1115*data_w +:data_w]), .r(v1115ibus), .q(v1115obus), .dec(dec[1115]));
wire [data_w*6-1:0] v1116ibus;
wire [temp_w*6-1:0] v1116obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1116 (.l(l[1116*data_w +:data_w]), .r(v1116ibus), .q(v1116obus), .dec(dec[1116]));
wire [data_w*6-1:0] v1117ibus;
wire [temp_w*6-1:0] v1117obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1117 (.l(l[1117*data_w +:data_w]), .r(v1117ibus), .q(v1117obus), .dec(dec[1117]));
wire [data_w*6-1:0] v1118ibus;
wire [temp_w*6-1:0] v1118obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1118 (.l(l[1118*data_w +:data_w]), .r(v1118ibus), .q(v1118obus), .dec(dec[1118]));
wire [data_w*6-1:0] v1119ibus;
wire [temp_w*6-1:0] v1119obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1119 (.l(l[1119*data_w +:data_w]), .r(v1119ibus), .q(v1119obus), .dec(dec[1119]));
wire [data_w*6-1:0] v1120ibus;
wire [temp_w*6-1:0] v1120obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1120 (.l(l[1120*data_w +:data_w]), .r(v1120ibus), .q(v1120obus), .dec(dec[1120]));
wire [data_w*6-1:0] v1121ibus;
wire [temp_w*6-1:0] v1121obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1121 (.l(l[1121*data_w +:data_w]), .r(v1121ibus), .q(v1121obus), .dec(dec[1121]));
wire [data_w*6-1:0] v1122ibus;
wire [temp_w*6-1:0] v1122obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1122 (.l(l[1122*data_w +:data_w]), .r(v1122ibus), .q(v1122obus), .dec(dec[1122]));
wire [data_w*6-1:0] v1123ibus;
wire [temp_w*6-1:0] v1123obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1123 (.l(l[1123*data_w +:data_w]), .r(v1123ibus), .q(v1123obus), .dec(dec[1123]));
wire [data_w*6-1:0] v1124ibus;
wire [temp_w*6-1:0] v1124obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1124 (.l(l[1124*data_w +:data_w]), .r(v1124ibus), .q(v1124obus), .dec(dec[1124]));
wire [data_w*6-1:0] v1125ibus;
wire [temp_w*6-1:0] v1125obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1125 (.l(l[1125*data_w +:data_w]), .r(v1125ibus), .q(v1125obus), .dec(dec[1125]));
wire [data_w*6-1:0] v1126ibus;
wire [temp_w*6-1:0] v1126obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1126 (.l(l[1126*data_w +:data_w]), .r(v1126ibus), .q(v1126obus), .dec(dec[1126]));
wire [data_w*6-1:0] v1127ibus;
wire [temp_w*6-1:0] v1127obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1127 (.l(l[1127*data_w +:data_w]), .r(v1127ibus), .q(v1127obus), .dec(dec[1127]));
wire [data_w*6-1:0] v1128ibus;
wire [temp_w*6-1:0] v1128obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1128 (.l(l[1128*data_w +:data_w]), .r(v1128ibus), .q(v1128obus), .dec(dec[1128]));
wire [data_w*6-1:0] v1129ibus;
wire [temp_w*6-1:0] v1129obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1129 (.l(l[1129*data_w +:data_w]), .r(v1129ibus), .q(v1129obus), .dec(dec[1129]));
wire [data_w*6-1:0] v1130ibus;
wire [temp_w*6-1:0] v1130obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1130 (.l(l[1130*data_w +:data_w]), .r(v1130ibus), .q(v1130obus), .dec(dec[1130]));
wire [data_w*6-1:0] v1131ibus;
wire [temp_w*6-1:0] v1131obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1131 (.l(l[1131*data_w +:data_w]), .r(v1131ibus), .q(v1131obus), .dec(dec[1131]));
wire [data_w*6-1:0] v1132ibus;
wire [temp_w*6-1:0] v1132obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1132 (.l(l[1132*data_w +:data_w]), .r(v1132ibus), .q(v1132obus), .dec(dec[1132]));
wire [data_w*6-1:0] v1133ibus;
wire [temp_w*6-1:0] v1133obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1133 (.l(l[1133*data_w +:data_w]), .r(v1133ibus), .q(v1133obus), .dec(dec[1133]));
wire [data_w*6-1:0] v1134ibus;
wire [temp_w*6-1:0] v1134obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1134 (.l(l[1134*data_w +:data_w]), .r(v1134ibus), .q(v1134obus), .dec(dec[1134]));
wire [data_w*6-1:0] v1135ibus;
wire [temp_w*6-1:0] v1135obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1135 (.l(l[1135*data_w +:data_w]), .r(v1135ibus), .q(v1135obus), .dec(dec[1135]));
wire [data_w*6-1:0] v1136ibus;
wire [temp_w*6-1:0] v1136obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1136 (.l(l[1136*data_w +:data_w]), .r(v1136ibus), .q(v1136obus), .dec(dec[1136]));
wire [data_w*6-1:0] v1137ibus;
wire [temp_w*6-1:0] v1137obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1137 (.l(l[1137*data_w +:data_w]), .r(v1137ibus), .q(v1137obus), .dec(dec[1137]));
wire [data_w*6-1:0] v1138ibus;
wire [temp_w*6-1:0] v1138obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1138 (.l(l[1138*data_w +:data_w]), .r(v1138ibus), .q(v1138obus), .dec(dec[1138]));
wire [data_w*6-1:0] v1139ibus;
wire [temp_w*6-1:0] v1139obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1139 (.l(l[1139*data_w +:data_w]), .r(v1139ibus), .q(v1139obus), .dec(dec[1139]));
wire [data_w*6-1:0] v1140ibus;
wire [temp_w*6-1:0] v1140obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1140 (.l(l[1140*data_w +:data_w]), .r(v1140ibus), .q(v1140obus), .dec(dec[1140]));
wire [data_w*6-1:0] v1141ibus;
wire [temp_w*6-1:0] v1141obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1141 (.l(l[1141*data_w +:data_w]), .r(v1141ibus), .q(v1141obus), .dec(dec[1141]));
wire [data_w*6-1:0] v1142ibus;
wire [temp_w*6-1:0] v1142obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1142 (.l(l[1142*data_w +:data_w]), .r(v1142ibus), .q(v1142obus), .dec(dec[1142]));
wire [data_w*6-1:0] v1143ibus;
wire [temp_w*6-1:0] v1143obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1143 (.l(l[1143*data_w +:data_w]), .r(v1143ibus), .q(v1143obus), .dec(dec[1143]));
wire [data_w*6-1:0] v1144ibus;
wire [temp_w*6-1:0] v1144obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1144 (.l(l[1144*data_w +:data_w]), .r(v1144ibus), .q(v1144obus), .dec(dec[1144]));
wire [data_w*6-1:0] v1145ibus;
wire [temp_w*6-1:0] v1145obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1145 (.l(l[1145*data_w +:data_w]), .r(v1145ibus), .q(v1145obus), .dec(dec[1145]));
wire [data_w*6-1:0] v1146ibus;
wire [temp_w*6-1:0] v1146obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1146 (.l(l[1146*data_w +:data_w]), .r(v1146ibus), .q(v1146obus), .dec(dec[1146]));
wire [data_w*6-1:0] v1147ibus;
wire [temp_w*6-1:0] v1147obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1147 (.l(l[1147*data_w +:data_w]), .r(v1147ibus), .q(v1147obus), .dec(dec[1147]));
wire [data_w*6-1:0] v1148ibus;
wire [temp_w*6-1:0] v1148obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1148 (.l(l[1148*data_w +:data_w]), .r(v1148ibus), .q(v1148obus), .dec(dec[1148]));
wire [data_w*6-1:0] v1149ibus;
wire [temp_w*6-1:0] v1149obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1149 (.l(l[1149*data_w +:data_w]), .r(v1149ibus), .q(v1149obus), .dec(dec[1149]));
wire [data_w*6-1:0] v1150ibus;
wire [temp_w*6-1:0] v1150obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1150 (.l(l[1150*data_w +:data_w]), .r(v1150ibus), .q(v1150obus), .dec(dec[1150]));
wire [data_w*6-1:0] v1151ibus;
wire [temp_w*6-1:0] v1151obus;
vnu #(.data_w(data_w), .D(6), .ext_w(ext_w)) VNU1151 (.l(l[1151*data_w +:data_w]), .r(v1151ibus), .q(v1151obus), .dec(dec[1151]));
wire [data_w*3-1:0] v1152ibus;
wire [temp_w*3-1:0] v1152obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1152 (.l(l[1152*data_w +:data_w]), .r(v1152ibus), .q(v1152obus), .dec(dec[1152]));
wire [data_w*3-1:0] v1153ibus;
wire [temp_w*3-1:0] v1153obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1153 (.l(l[1153*data_w +:data_w]), .r(v1153ibus), .q(v1153obus), .dec(dec[1153]));
wire [data_w*3-1:0] v1154ibus;
wire [temp_w*3-1:0] v1154obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1154 (.l(l[1154*data_w +:data_w]), .r(v1154ibus), .q(v1154obus), .dec(dec[1154]));
wire [data_w*3-1:0] v1155ibus;
wire [temp_w*3-1:0] v1155obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1155 (.l(l[1155*data_w +:data_w]), .r(v1155ibus), .q(v1155obus), .dec(dec[1155]));
wire [data_w*3-1:0] v1156ibus;
wire [temp_w*3-1:0] v1156obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1156 (.l(l[1156*data_w +:data_w]), .r(v1156ibus), .q(v1156obus), .dec(dec[1156]));
wire [data_w*3-1:0] v1157ibus;
wire [temp_w*3-1:0] v1157obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1157 (.l(l[1157*data_w +:data_w]), .r(v1157ibus), .q(v1157obus), .dec(dec[1157]));
wire [data_w*3-1:0] v1158ibus;
wire [temp_w*3-1:0] v1158obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1158 (.l(l[1158*data_w +:data_w]), .r(v1158ibus), .q(v1158obus), .dec(dec[1158]));
wire [data_w*3-1:0] v1159ibus;
wire [temp_w*3-1:0] v1159obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1159 (.l(l[1159*data_w +:data_w]), .r(v1159ibus), .q(v1159obus), .dec(dec[1159]));
wire [data_w*3-1:0] v1160ibus;
wire [temp_w*3-1:0] v1160obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1160 (.l(l[1160*data_w +:data_w]), .r(v1160ibus), .q(v1160obus), .dec(dec[1160]));
wire [data_w*3-1:0] v1161ibus;
wire [temp_w*3-1:0] v1161obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1161 (.l(l[1161*data_w +:data_w]), .r(v1161ibus), .q(v1161obus), .dec(dec[1161]));
wire [data_w*3-1:0] v1162ibus;
wire [temp_w*3-1:0] v1162obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1162 (.l(l[1162*data_w +:data_w]), .r(v1162ibus), .q(v1162obus), .dec(dec[1162]));
wire [data_w*3-1:0] v1163ibus;
wire [temp_w*3-1:0] v1163obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1163 (.l(l[1163*data_w +:data_w]), .r(v1163ibus), .q(v1163obus), .dec(dec[1163]));
wire [data_w*3-1:0] v1164ibus;
wire [temp_w*3-1:0] v1164obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1164 (.l(l[1164*data_w +:data_w]), .r(v1164ibus), .q(v1164obus), .dec(dec[1164]));
wire [data_w*3-1:0] v1165ibus;
wire [temp_w*3-1:0] v1165obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1165 (.l(l[1165*data_w +:data_w]), .r(v1165ibus), .q(v1165obus), .dec(dec[1165]));
wire [data_w*3-1:0] v1166ibus;
wire [temp_w*3-1:0] v1166obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1166 (.l(l[1166*data_w +:data_w]), .r(v1166ibus), .q(v1166obus), .dec(dec[1166]));
wire [data_w*3-1:0] v1167ibus;
wire [temp_w*3-1:0] v1167obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1167 (.l(l[1167*data_w +:data_w]), .r(v1167ibus), .q(v1167obus), .dec(dec[1167]));
wire [data_w*3-1:0] v1168ibus;
wire [temp_w*3-1:0] v1168obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1168 (.l(l[1168*data_w +:data_w]), .r(v1168ibus), .q(v1168obus), .dec(dec[1168]));
wire [data_w*3-1:0] v1169ibus;
wire [temp_w*3-1:0] v1169obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1169 (.l(l[1169*data_w +:data_w]), .r(v1169ibus), .q(v1169obus), .dec(dec[1169]));
wire [data_w*3-1:0] v1170ibus;
wire [temp_w*3-1:0] v1170obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1170 (.l(l[1170*data_w +:data_w]), .r(v1170ibus), .q(v1170obus), .dec(dec[1170]));
wire [data_w*3-1:0] v1171ibus;
wire [temp_w*3-1:0] v1171obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1171 (.l(l[1171*data_w +:data_w]), .r(v1171ibus), .q(v1171obus), .dec(dec[1171]));
wire [data_w*3-1:0] v1172ibus;
wire [temp_w*3-1:0] v1172obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1172 (.l(l[1172*data_w +:data_w]), .r(v1172ibus), .q(v1172obus), .dec(dec[1172]));
wire [data_w*3-1:0] v1173ibus;
wire [temp_w*3-1:0] v1173obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1173 (.l(l[1173*data_w +:data_w]), .r(v1173ibus), .q(v1173obus), .dec(dec[1173]));
wire [data_w*3-1:0] v1174ibus;
wire [temp_w*3-1:0] v1174obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1174 (.l(l[1174*data_w +:data_w]), .r(v1174ibus), .q(v1174obus), .dec(dec[1174]));
wire [data_w*3-1:0] v1175ibus;
wire [temp_w*3-1:0] v1175obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1175 (.l(l[1175*data_w +:data_w]), .r(v1175ibus), .q(v1175obus), .dec(dec[1175]));
wire [data_w*3-1:0] v1176ibus;
wire [temp_w*3-1:0] v1176obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1176 (.l(l[1176*data_w +:data_w]), .r(v1176ibus), .q(v1176obus), .dec(dec[1176]));
wire [data_w*3-1:0] v1177ibus;
wire [temp_w*3-1:0] v1177obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1177 (.l(l[1177*data_w +:data_w]), .r(v1177ibus), .q(v1177obus), .dec(dec[1177]));
wire [data_w*3-1:0] v1178ibus;
wire [temp_w*3-1:0] v1178obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1178 (.l(l[1178*data_w +:data_w]), .r(v1178ibus), .q(v1178obus), .dec(dec[1178]));
wire [data_w*3-1:0] v1179ibus;
wire [temp_w*3-1:0] v1179obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1179 (.l(l[1179*data_w +:data_w]), .r(v1179ibus), .q(v1179obus), .dec(dec[1179]));
wire [data_w*3-1:0] v1180ibus;
wire [temp_w*3-1:0] v1180obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1180 (.l(l[1180*data_w +:data_w]), .r(v1180ibus), .q(v1180obus), .dec(dec[1180]));
wire [data_w*3-1:0] v1181ibus;
wire [temp_w*3-1:0] v1181obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1181 (.l(l[1181*data_w +:data_w]), .r(v1181ibus), .q(v1181obus), .dec(dec[1181]));
wire [data_w*3-1:0] v1182ibus;
wire [temp_w*3-1:0] v1182obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1182 (.l(l[1182*data_w +:data_w]), .r(v1182ibus), .q(v1182obus), .dec(dec[1182]));
wire [data_w*3-1:0] v1183ibus;
wire [temp_w*3-1:0] v1183obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1183 (.l(l[1183*data_w +:data_w]), .r(v1183ibus), .q(v1183obus), .dec(dec[1183]));
wire [data_w*3-1:0] v1184ibus;
wire [temp_w*3-1:0] v1184obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1184 (.l(l[1184*data_w +:data_w]), .r(v1184ibus), .q(v1184obus), .dec(dec[1184]));
wire [data_w*3-1:0] v1185ibus;
wire [temp_w*3-1:0] v1185obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1185 (.l(l[1185*data_w +:data_w]), .r(v1185ibus), .q(v1185obus), .dec(dec[1185]));
wire [data_w*3-1:0] v1186ibus;
wire [temp_w*3-1:0] v1186obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1186 (.l(l[1186*data_w +:data_w]), .r(v1186ibus), .q(v1186obus), .dec(dec[1186]));
wire [data_w*3-1:0] v1187ibus;
wire [temp_w*3-1:0] v1187obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1187 (.l(l[1187*data_w +:data_w]), .r(v1187ibus), .q(v1187obus), .dec(dec[1187]));
wire [data_w*3-1:0] v1188ibus;
wire [temp_w*3-1:0] v1188obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1188 (.l(l[1188*data_w +:data_w]), .r(v1188ibus), .q(v1188obus), .dec(dec[1188]));
wire [data_w*3-1:0] v1189ibus;
wire [temp_w*3-1:0] v1189obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1189 (.l(l[1189*data_w +:data_w]), .r(v1189ibus), .q(v1189obus), .dec(dec[1189]));
wire [data_w*3-1:0] v1190ibus;
wire [temp_w*3-1:0] v1190obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1190 (.l(l[1190*data_w +:data_w]), .r(v1190ibus), .q(v1190obus), .dec(dec[1190]));
wire [data_w*3-1:0] v1191ibus;
wire [temp_w*3-1:0] v1191obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1191 (.l(l[1191*data_w +:data_w]), .r(v1191ibus), .q(v1191obus), .dec(dec[1191]));
wire [data_w*3-1:0] v1192ibus;
wire [temp_w*3-1:0] v1192obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1192 (.l(l[1192*data_w +:data_w]), .r(v1192ibus), .q(v1192obus), .dec(dec[1192]));
wire [data_w*3-1:0] v1193ibus;
wire [temp_w*3-1:0] v1193obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1193 (.l(l[1193*data_w +:data_w]), .r(v1193ibus), .q(v1193obus), .dec(dec[1193]));
wire [data_w*3-1:0] v1194ibus;
wire [temp_w*3-1:0] v1194obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1194 (.l(l[1194*data_w +:data_w]), .r(v1194ibus), .q(v1194obus), .dec(dec[1194]));
wire [data_w*3-1:0] v1195ibus;
wire [temp_w*3-1:0] v1195obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1195 (.l(l[1195*data_w +:data_w]), .r(v1195ibus), .q(v1195obus), .dec(dec[1195]));
wire [data_w*3-1:0] v1196ibus;
wire [temp_w*3-1:0] v1196obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1196 (.l(l[1196*data_w +:data_w]), .r(v1196ibus), .q(v1196obus), .dec(dec[1196]));
wire [data_w*3-1:0] v1197ibus;
wire [temp_w*3-1:0] v1197obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1197 (.l(l[1197*data_w +:data_w]), .r(v1197ibus), .q(v1197obus), .dec(dec[1197]));
wire [data_w*3-1:0] v1198ibus;
wire [temp_w*3-1:0] v1198obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1198 (.l(l[1198*data_w +:data_w]), .r(v1198ibus), .q(v1198obus), .dec(dec[1198]));
wire [data_w*3-1:0] v1199ibus;
wire [temp_w*3-1:0] v1199obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1199 (.l(l[1199*data_w +:data_w]), .r(v1199ibus), .q(v1199obus), .dec(dec[1199]));
wire [data_w*3-1:0] v1200ibus;
wire [temp_w*3-1:0] v1200obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1200 (.l(l[1200*data_w +:data_w]), .r(v1200ibus), .q(v1200obus), .dec(dec[1200]));
wire [data_w*3-1:0] v1201ibus;
wire [temp_w*3-1:0] v1201obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1201 (.l(l[1201*data_w +:data_w]), .r(v1201ibus), .q(v1201obus), .dec(dec[1201]));
wire [data_w*3-1:0] v1202ibus;
wire [temp_w*3-1:0] v1202obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1202 (.l(l[1202*data_w +:data_w]), .r(v1202ibus), .q(v1202obus), .dec(dec[1202]));
wire [data_w*3-1:0] v1203ibus;
wire [temp_w*3-1:0] v1203obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1203 (.l(l[1203*data_w +:data_w]), .r(v1203ibus), .q(v1203obus), .dec(dec[1203]));
wire [data_w*3-1:0] v1204ibus;
wire [temp_w*3-1:0] v1204obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1204 (.l(l[1204*data_w +:data_w]), .r(v1204ibus), .q(v1204obus), .dec(dec[1204]));
wire [data_w*3-1:0] v1205ibus;
wire [temp_w*3-1:0] v1205obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1205 (.l(l[1205*data_w +:data_w]), .r(v1205ibus), .q(v1205obus), .dec(dec[1205]));
wire [data_w*3-1:0] v1206ibus;
wire [temp_w*3-1:0] v1206obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1206 (.l(l[1206*data_w +:data_w]), .r(v1206ibus), .q(v1206obus), .dec(dec[1206]));
wire [data_w*3-1:0] v1207ibus;
wire [temp_w*3-1:0] v1207obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1207 (.l(l[1207*data_w +:data_w]), .r(v1207ibus), .q(v1207obus), .dec(dec[1207]));
wire [data_w*3-1:0] v1208ibus;
wire [temp_w*3-1:0] v1208obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1208 (.l(l[1208*data_w +:data_w]), .r(v1208ibus), .q(v1208obus), .dec(dec[1208]));
wire [data_w*3-1:0] v1209ibus;
wire [temp_w*3-1:0] v1209obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1209 (.l(l[1209*data_w +:data_w]), .r(v1209ibus), .q(v1209obus), .dec(dec[1209]));
wire [data_w*3-1:0] v1210ibus;
wire [temp_w*3-1:0] v1210obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1210 (.l(l[1210*data_w +:data_w]), .r(v1210ibus), .q(v1210obus), .dec(dec[1210]));
wire [data_w*3-1:0] v1211ibus;
wire [temp_w*3-1:0] v1211obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1211 (.l(l[1211*data_w +:data_w]), .r(v1211ibus), .q(v1211obus), .dec(dec[1211]));
wire [data_w*3-1:0] v1212ibus;
wire [temp_w*3-1:0] v1212obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1212 (.l(l[1212*data_w +:data_w]), .r(v1212ibus), .q(v1212obus), .dec(dec[1212]));
wire [data_w*3-1:0] v1213ibus;
wire [temp_w*3-1:0] v1213obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1213 (.l(l[1213*data_w +:data_w]), .r(v1213ibus), .q(v1213obus), .dec(dec[1213]));
wire [data_w*3-1:0] v1214ibus;
wire [temp_w*3-1:0] v1214obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1214 (.l(l[1214*data_w +:data_w]), .r(v1214ibus), .q(v1214obus), .dec(dec[1214]));
wire [data_w*3-1:0] v1215ibus;
wire [temp_w*3-1:0] v1215obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1215 (.l(l[1215*data_w +:data_w]), .r(v1215ibus), .q(v1215obus), .dec(dec[1215]));
wire [data_w*3-1:0] v1216ibus;
wire [temp_w*3-1:0] v1216obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1216 (.l(l[1216*data_w +:data_w]), .r(v1216ibus), .q(v1216obus), .dec(dec[1216]));
wire [data_w*3-1:0] v1217ibus;
wire [temp_w*3-1:0] v1217obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1217 (.l(l[1217*data_w +:data_w]), .r(v1217ibus), .q(v1217obus), .dec(dec[1217]));
wire [data_w*3-1:0] v1218ibus;
wire [temp_w*3-1:0] v1218obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1218 (.l(l[1218*data_w +:data_w]), .r(v1218ibus), .q(v1218obus), .dec(dec[1218]));
wire [data_w*3-1:0] v1219ibus;
wire [temp_w*3-1:0] v1219obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1219 (.l(l[1219*data_w +:data_w]), .r(v1219ibus), .q(v1219obus), .dec(dec[1219]));
wire [data_w*3-1:0] v1220ibus;
wire [temp_w*3-1:0] v1220obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1220 (.l(l[1220*data_w +:data_w]), .r(v1220ibus), .q(v1220obus), .dec(dec[1220]));
wire [data_w*3-1:0] v1221ibus;
wire [temp_w*3-1:0] v1221obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1221 (.l(l[1221*data_w +:data_w]), .r(v1221ibus), .q(v1221obus), .dec(dec[1221]));
wire [data_w*3-1:0] v1222ibus;
wire [temp_w*3-1:0] v1222obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1222 (.l(l[1222*data_w +:data_w]), .r(v1222ibus), .q(v1222obus), .dec(dec[1222]));
wire [data_w*3-1:0] v1223ibus;
wire [temp_w*3-1:0] v1223obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1223 (.l(l[1223*data_w +:data_w]), .r(v1223ibus), .q(v1223obus), .dec(dec[1223]));
wire [data_w*3-1:0] v1224ibus;
wire [temp_w*3-1:0] v1224obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1224 (.l(l[1224*data_w +:data_w]), .r(v1224ibus), .q(v1224obus), .dec(dec[1224]));
wire [data_w*3-1:0] v1225ibus;
wire [temp_w*3-1:0] v1225obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1225 (.l(l[1225*data_w +:data_w]), .r(v1225ibus), .q(v1225obus), .dec(dec[1225]));
wire [data_w*3-1:0] v1226ibus;
wire [temp_w*3-1:0] v1226obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1226 (.l(l[1226*data_w +:data_w]), .r(v1226ibus), .q(v1226obus), .dec(dec[1226]));
wire [data_w*3-1:0] v1227ibus;
wire [temp_w*3-1:0] v1227obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1227 (.l(l[1227*data_w +:data_w]), .r(v1227ibus), .q(v1227obus), .dec(dec[1227]));
wire [data_w*3-1:0] v1228ibus;
wire [temp_w*3-1:0] v1228obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1228 (.l(l[1228*data_w +:data_w]), .r(v1228ibus), .q(v1228obus), .dec(dec[1228]));
wire [data_w*3-1:0] v1229ibus;
wire [temp_w*3-1:0] v1229obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1229 (.l(l[1229*data_w +:data_w]), .r(v1229ibus), .q(v1229obus), .dec(dec[1229]));
wire [data_w*3-1:0] v1230ibus;
wire [temp_w*3-1:0] v1230obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1230 (.l(l[1230*data_w +:data_w]), .r(v1230ibus), .q(v1230obus), .dec(dec[1230]));
wire [data_w*3-1:0] v1231ibus;
wire [temp_w*3-1:0] v1231obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1231 (.l(l[1231*data_w +:data_w]), .r(v1231ibus), .q(v1231obus), .dec(dec[1231]));
wire [data_w*3-1:0] v1232ibus;
wire [temp_w*3-1:0] v1232obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1232 (.l(l[1232*data_w +:data_w]), .r(v1232ibus), .q(v1232obus), .dec(dec[1232]));
wire [data_w*3-1:0] v1233ibus;
wire [temp_w*3-1:0] v1233obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1233 (.l(l[1233*data_w +:data_w]), .r(v1233ibus), .q(v1233obus), .dec(dec[1233]));
wire [data_w*3-1:0] v1234ibus;
wire [temp_w*3-1:0] v1234obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1234 (.l(l[1234*data_w +:data_w]), .r(v1234ibus), .q(v1234obus), .dec(dec[1234]));
wire [data_w*3-1:0] v1235ibus;
wire [temp_w*3-1:0] v1235obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1235 (.l(l[1235*data_w +:data_w]), .r(v1235ibus), .q(v1235obus), .dec(dec[1235]));
wire [data_w*3-1:0] v1236ibus;
wire [temp_w*3-1:0] v1236obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1236 (.l(l[1236*data_w +:data_w]), .r(v1236ibus), .q(v1236obus), .dec(dec[1236]));
wire [data_w*3-1:0] v1237ibus;
wire [temp_w*3-1:0] v1237obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1237 (.l(l[1237*data_w +:data_w]), .r(v1237ibus), .q(v1237obus), .dec(dec[1237]));
wire [data_w*3-1:0] v1238ibus;
wire [temp_w*3-1:0] v1238obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1238 (.l(l[1238*data_w +:data_w]), .r(v1238ibus), .q(v1238obus), .dec(dec[1238]));
wire [data_w*3-1:0] v1239ibus;
wire [temp_w*3-1:0] v1239obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1239 (.l(l[1239*data_w +:data_w]), .r(v1239ibus), .q(v1239obus), .dec(dec[1239]));
wire [data_w*3-1:0] v1240ibus;
wire [temp_w*3-1:0] v1240obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1240 (.l(l[1240*data_w +:data_w]), .r(v1240ibus), .q(v1240obus), .dec(dec[1240]));
wire [data_w*3-1:0] v1241ibus;
wire [temp_w*3-1:0] v1241obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1241 (.l(l[1241*data_w +:data_w]), .r(v1241ibus), .q(v1241obus), .dec(dec[1241]));
wire [data_w*3-1:0] v1242ibus;
wire [temp_w*3-1:0] v1242obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1242 (.l(l[1242*data_w +:data_w]), .r(v1242ibus), .q(v1242obus), .dec(dec[1242]));
wire [data_w*3-1:0] v1243ibus;
wire [temp_w*3-1:0] v1243obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1243 (.l(l[1243*data_w +:data_w]), .r(v1243ibus), .q(v1243obus), .dec(dec[1243]));
wire [data_w*3-1:0] v1244ibus;
wire [temp_w*3-1:0] v1244obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1244 (.l(l[1244*data_w +:data_w]), .r(v1244ibus), .q(v1244obus), .dec(dec[1244]));
wire [data_w*3-1:0] v1245ibus;
wire [temp_w*3-1:0] v1245obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1245 (.l(l[1245*data_w +:data_w]), .r(v1245ibus), .q(v1245obus), .dec(dec[1245]));
wire [data_w*3-1:0] v1246ibus;
wire [temp_w*3-1:0] v1246obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1246 (.l(l[1246*data_w +:data_w]), .r(v1246ibus), .q(v1246obus), .dec(dec[1246]));
wire [data_w*3-1:0] v1247ibus;
wire [temp_w*3-1:0] v1247obus;
vnu #(.data_w(data_w), .D(3), .ext_w(ext_w)) VNU1247 (.l(l[1247*data_w +:data_w]), .r(v1247ibus), .q(v1247obus), .dec(dec[1247]));
wire [data_w*2-1:0] v1248ibus;
wire [temp_w*2-1:0] v1248obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1248 (.l(l[1248*data_w +:data_w]), .r(v1248ibus), .q(v1248obus), .dec(dec[1248]));
wire [data_w*2-1:0] v1249ibus;
wire [temp_w*2-1:0] v1249obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1249 (.l(l[1249*data_w +:data_w]), .r(v1249ibus), .q(v1249obus), .dec(dec[1249]));
wire [data_w*2-1:0] v1250ibus;
wire [temp_w*2-1:0] v1250obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1250 (.l(l[1250*data_w +:data_w]), .r(v1250ibus), .q(v1250obus), .dec(dec[1250]));
wire [data_w*2-1:0] v1251ibus;
wire [temp_w*2-1:0] v1251obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1251 (.l(l[1251*data_w +:data_w]), .r(v1251ibus), .q(v1251obus), .dec(dec[1251]));
wire [data_w*2-1:0] v1252ibus;
wire [temp_w*2-1:0] v1252obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1252 (.l(l[1252*data_w +:data_w]), .r(v1252ibus), .q(v1252obus), .dec(dec[1252]));
wire [data_w*2-1:0] v1253ibus;
wire [temp_w*2-1:0] v1253obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1253 (.l(l[1253*data_w +:data_w]), .r(v1253ibus), .q(v1253obus), .dec(dec[1253]));
wire [data_w*2-1:0] v1254ibus;
wire [temp_w*2-1:0] v1254obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1254 (.l(l[1254*data_w +:data_w]), .r(v1254ibus), .q(v1254obus), .dec(dec[1254]));
wire [data_w*2-1:0] v1255ibus;
wire [temp_w*2-1:0] v1255obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1255 (.l(l[1255*data_w +:data_w]), .r(v1255ibus), .q(v1255obus), .dec(dec[1255]));
wire [data_w*2-1:0] v1256ibus;
wire [temp_w*2-1:0] v1256obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1256 (.l(l[1256*data_w +:data_w]), .r(v1256ibus), .q(v1256obus), .dec(dec[1256]));
wire [data_w*2-1:0] v1257ibus;
wire [temp_w*2-1:0] v1257obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1257 (.l(l[1257*data_w +:data_w]), .r(v1257ibus), .q(v1257obus), .dec(dec[1257]));
wire [data_w*2-1:0] v1258ibus;
wire [temp_w*2-1:0] v1258obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1258 (.l(l[1258*data_w +:data_w]), .r(v1258ibus), .q(v1258obus), .dec(dec[1258]));
wire [data_w*2-1:0] v1259ibus;
wire [temp_w*2-1:0] v1259obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1259 (.l(l[1259*data_w +:data_w]), .r(v1259ibus), .q(v1259obus), .dec(dec[1259]));
wire [data_w*2-1:0] v1260ibus;
wire [temp_w*2-1:0] v1260obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1260 (.l(l[1260*data_w +:data_w]), .r(v1260ibus), .q(v1260obus), .dec(dec[1260]));
wire [data_w*2-1:0] v1261ibus;
wire [temp_w*2-1:0] v1261obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1261 (.l(l[1261*data_w +:data_w]), .r(v1261ibus), .q(v1261obus), .dec(dec[1261]));
wire [data_w*2-1:0] v1262ibus;
wire [temp_w*2-1:0] v1262obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1262 (.l(l[1262*data_w +:data_w]), .r(v1262ibus), .q(v1262obus), .dec(dec[1262]));
wire [data_w*2-1:0] v1263ibus;
wire [temp_w*2-1:0] v1263obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1263 (.l(l[1263*data_w +:data_w]), .r(v1263ibus), .q(v1263obus), .dec(dec[1263]));
wire [data_w*2-1:0] v1264ibus;
wire [temp_w*2-1:0] v1264obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1264 (.l(l[1264*data_w +:data_w]), .r(v1264ibus), .q(v1264obus), .dec(dec[1264]));
wire [data_w*2-1:0] v1265ibus;
wire [temp_w*2-1:0] v1265obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1265 (.l(l[1265*data_w +:data_w]), .r(v1265ibus), .q(v1265obus), .dec(dec[1265]));
wire [data_w*2-1:0] v1266ibus;
wire [temp_w*2-1:0] v1266obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1266 (.l(l[1266*data_w +:data_w]), .r(v1266ibus), .q(v1266obus), .dec(dec[1266]));
wire [data_w*2-1:0] v1267ibus;
wire [temp_w*2-1:0] v1267obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1267 (.l(l[1267*data_w +:data_w]), .r(v1267ibus), .q(v1267obus), .dec(dec[1267]));
wire [data_w*2-1:0] v1268ibus;
wire [temp_w*2-1:0] v1268obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1268 (.l(l[1268*data_w +:data_w]), .r(v1268ibus), .q(v1268obus), .dec(dec[1268]));
wire [data_w*2-1:0] v1269ibus;
wire [temp_w*2-1:0] v1269obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1269 (.l(l[1269*data_w +:data_w]), .r(v1269ibus), .q(v1269obus), .dec(dec[1269]));
wire [data_w*2-1:0] v1270ibus;
wire [temp_w*2-1:0] v1270obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1270 (.l(l[1270*data_w +:data_w]), .r(v1270ibus), .q(v1270obus), .dec(dec[1270]));
wire [data_w*2-1:0] v1271ibus;
wire [temp_w*2-1:0] v1271obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1271 (.l(l[1271*data_w +:data_w]), .r(v1271ibus), .q(v1271obus), .dec(dec[1271]));
wire [data_w*2-1:0] v1272ibus;
wire [temp_w*2-1:0] v1272obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1272 (.l(l[1272*data_w +:data_w]), .r(v1272ibus), .q(v1272obus), .dec(dec[1272]));
wire [data_w*2-1:0] v1273ibus;
wire [temp_w*2-1:0] v1273obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1273 (.l(l[1273*data_w +:data_w]), .r(v1273ibus), .q(v1273obus), .dec(dec[1273]));
wire [data_w*2-1:0] v1274ibus;
wire [temp_w*2-1:0] v1274obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1274 (.l(l[1274*data_w +:data_w]), .r(v1274ibus), .q(v1274obus), .dec(dec[1274]));
wire [data_w*2-1:0] v1275ibus;
wire [temp_w*2-1:0] v1275obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1275 (.l(l[1275*data_w +:data_w]), .r(v1275ibus), .q(v1275obus), .dec(dec[1275]));
wire [data_w*2-1:0] v1276ibus;
wire [temp_w*2-1:0] v1276obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1276 (.l(l[1276*data_w +:data_w]), .r(v1276ibus), .q(v1276obus), .dec(dec[1276]));
wire [data_w*2-1:0] v1277ibus;
wire [temp_w*2-1:0] v1277obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1277 (.l(l[1277*data_w +:data_w]), .r(v1277ibus), .q(v1277obus), .dec(dec[1277]));
wire [data_w*2-1:0] v1278ibus;
wire [temp_w*2-1:0] v1278obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1278 (.l(l[1278*data_w +:data_w]), .r(v1278ibus), .q(v1278obus), .dec(dec[1278]));
wire [data_w*2-1:0] v1279ibus;
wire [temp_w*2-1:0] v1279obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1279 (.l(l[1279*data_w +:data_w]), .r(v1279ibus), .q(v1279obus), .dec(dec[1279]));
wire [data_w*2-1:0] v1280ibus;
wire [temp_w*2-1:0] v1280obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1280 (.l(l[1280*data_w +:data_w]), .r(v1280ibus), .q(v1280obus), .dec(dec[1280]));
wire [data_w*2-1:0] v1281ibus;
wire [temp_w*2-1:0] v1281obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1281 (.l(l[1281*data_w +:data_w]), .r(v1281ibus), .q(v1281obus), .dec(dec[1281]));
wire [data_w*2-1:0] v1282ibus;
wire [temp_w*2-1:0] v1282obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1282 (.l(l[1282*data_w +:data_w]), .r(v1282ibus), .q(v1282obus), .dec(dec[1282]));
wire [data_w*2-1:0] v1283ibus;
wire [temp_w*2-1:0] v1283obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1283 (.l(l[1283*data_w +:data_w]), .r(v1283ibus), .q(v1283obus), .dec(dec[1283]));
wire [data_w*2-1:0] v1284ibus;
wire [temp_w*2-1:0] v1284obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1284 (.l(l[1284*data_w +:data_w]), .r(v1284ibus), .q(v1284obus), .dec(dec[1284]));
wire [data_w*2-1:0] v1285ibus;
wire [temp_w*2-1:0] v1285obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1285 (.l(l[1285*data_w +:data_w]), .r(v1285ibus), .q(v1285obus), .dec(dec[1285]));
wire [data_w*2-1:0] v1286ibus;
wire [temp_w*2-1:0] v1286obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1286 (.l(l[1286*data_w +:data_w]), .r(v1286ibus), .q(v1286obus), .dec(dec[1286]));
wire [data_w*2-1:0] v1287ibus;
wire [temp_w*2-1:0] v1287obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1287 (.l(l[1287*data_w +:data_w]), .r(v1287ibus), .q(v1287obus), .dec(dec[1287]));
wire [data_w*2-1:0] v1288ibus;
wire [temp_w*2-1:0] v1288obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1288 (.l(l[1288*data_w +:data_w]), .r(v1288ibus), .q(v1288obus), .dec(dec[1288]));
wire [data_w*2-1:0] v1289ibus;
wire [temp_w*2-1:0] v1289obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1289 (.l(l[1289*data_w +:data_w]), .r(v1289ibus), .q(v1289obus), .dec(dec[1289]));
wire [data_w*2-1:0] v1290ibus;
wire [temp_w*2-1:0] v1290obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1290 (.l(l[1290*data_w +:data_w]), .r(v1290ibus), .q(v1290obus), .dec(dec[1290]));
wire [data_w*2-1:0] v1291ibus;
wire [temp_w*2-1:0] v1291obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1291 (.l(l[1291*data_w +:data_w]), .r(v1291ibus), .q(v1291obus), .dec(dec[1291]));
wire [data_w*2-1:0] v1292ibus;
wire [temp_w*2-1:0] v1292obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1292 (.l(l[1292*data_w +:data_w]), .r(v1292ibus), .q(v1292obus), .dec(dec[1292]));
wire [data_w*2-1:0] v1293ibus;
wire [temp_w*2-1:0] v1293obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1293 (.l(l[1293*data_w +:data_w]), .r(v1293ibus), .q(v1293obus), .dec(dec[1293]));
wire [data_w*2-1:0] v1294ibus;
wire [temp_w*2-1:0] v1294obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1294 (.l(l[1294*data_w +:data_w]), .r(v1294ibus), .q(v1294obus), .dec(dec[1294]));
wire [data_w*2-1:0] v1295ibus;
wire [temp_w*2-1:0] v1295obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1295 (.l(l[1295*data_w +:data_w]), .r(v1295ibus), .q(v1295obus), .dec(dec[1295]));
wire [data_w*2-1:0] v1296ibus;
wire [temp_w*2-1:0] v1296obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1296 (.l(l[1296*data_w +:data_w]), .r(v1296ibus), .q(v1296obus), .dec(dec[1296]));
wire [data_w*2-1:0] v1297ibus;
wire [temp_w*2-1:0] v1297obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1297 (.l(l[1297*data_w +:data_w]), .r(v1297ibus), .q(v1297obus), .dec(dec[1297]));
wire [data_w*2-1:0] v1298ibus;
wire [temp_w*2-1:0] v1298obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1298 (.l(l[1298*data_w +:data_w]), .r(v1298ibus), .q(v1298obus), .dec(dec[1298]));
wire [data_w*2-1:0] v1299ibus;
wire [temp_w*2-1:0] v1299obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1299 (.l(l[1299*data_w +:data_w]), .r(v1299ibus), .q(v1299obus), .dec(dec[1299]));
wire [data_w*2-1:0] v1300ibus;
wire [temp_w*2-1:0] v1300obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1300 (.l(l[1300*data_w +:data_w]), .r(v1300ibus), .q(v1300obus), .dec(dec[1300]));
wire [data_w*2-1:0] v1301ibus;
wire [temp_w*2-1:0] v1301obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1301 (.l(l[1301*data_w +:data_w]), .r(v1301ibus), .q(v1301obus), .dec(dec[1301]));
wire [data_w*2-1:0] v1302ibus;
wire [temp_w*2-1:0] v1302obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1302 (.l(l[1302*data_w +:data_w]), .r(v1302ibus), .q(v1302obus), .dec(dec[1302]));
wire [data_w*2-1:0] v1303ibus;
wire [temp_w*2-1:0] v1303obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1303 (.l(l[1303*data_w +:data_w]), .r(v1303ibus), .q(v1303obus), .dec(dec[1303]));
wire [data_w*2-1:0] v1304ibus;
wire [temp_w*2-1:0] v1304obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1304 (.l(l[1304*data_w +:data_w]), .r(v1304ibus), .q(v1304obus), .dec(dec[1304]));
wire [data_w*2-1:0] v1305ibus;
wire [temp_w*2-1:0] v1305obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1305 (.l(l[1305*data_w +:data_w]), .r(v1305ibus), .q(v1305obus), .dec(dec[1305]));
wire [data_w*2-1:0] v1306ibus;
wire [temp_w*2-1:0] v1306obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1306 (.l(l[1306*data_w +:data_w]), .r(v1306ibus), .q(v1306obus), .dec(dec[1306]));
wire [data_w*2-1:0] v1307ibus;
wire [temp_w*2-1:0] v1307obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1307 (.l(l[1307*data_w +:data_w]), .r(v1307ibus), .q(v1307obus), .dec(dec[1307]));
wire [data_w*2-1:0] v1308ibus;
wire [temp_w*2-1:0] v1308obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1308 (.l(l[1308*data_w +:data_w]), .r(v1308ibus), .q(v1308obus), .dec(dec[1308]));
wire [data_w*2-1:0] v1309ibus;
wire [temp_w*2-1:0] v1309obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1309 (.l(l[1309*data_w +:data_w]), .r(v1309ibus), .q(v1309obus), .dec(dec[1309]));
wire [data_w*2-1:0] v1310ibus;
wire [temp_w*2-1:0] v1310obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1310 (.l(l[1310*data_w +:data_w]), .r(v1310ibus), .q(v1310obus), .dec(dec[1310]));
wire [data_w*2-1:0] v1311ibus;
wire [temp_w*2-1:0] v1311obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1311 (.l(l[1311*data_w +:data_w]), .r(v1311ibus), .q(v1311obus), .dec(dec[1311]));
wire [data_w*2-1:0] v1312ibus;
wire [temp_w*2-1:0] v1312obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1312 (.l(l[1312*data_w +:data_w]), .r(v1312ibus), .q(v1312obus), .dec(dec[1312]));
wire [data_w*2-1:0] v1313ibus;
wire [temp_w*2-1:0] v1313obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1313 (.l(l[1313*data_w +:data_w]), .r(v1313ibus), .q(v1313obus), .dec(dec[1313]));
wire [data_w*2-1:0] v1314ibus;
wire [temp_w*2-1:0] v1314obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1314 (.l(l[1314*data_w +:data_w]), .r(v1314ibus), .q(v1314obus), .dec(dec[1314]));
wire [data_w*2-1:0] v1315ibus;
wire [temp_w*2-1:0] v1315obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1315 (.l(l[1315*data_w +:data_w]), .r(v1315ibus), .q(v1315obus), .dec(dec[1315]));
wire [data_w*2-1:0] v1316ibus;
wire [temp_w*2-1:0] v1316obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1316 (.l(l[1316*data_w +:data_w]), .r(v1316ibus), .q(v1316obus), .dec(dec[1316]));
wire [data_w*2-1:0] v1317ibus;
wire [temp_w*2-1:0] v1317obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1317 (.l(l[1317*data_w +:data_w]), .r(v1317ibus), .q(v1317obus), .dec(dec[1317]));
wire [data_w*2-1:0] v1318ibus;
wire [temp_w*2-1:0] v1318obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1318 (.l(l[1318*data_w +:data_w]), .r(v1318ibus), .q(v1318obus), .dec(dec[1318]));
wire [data_w*2-1:0] v1319ibus;
wire [temp_w*2-1:0] v1319obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1319 (.l(l[1319*data_w +:data_w]), .r(v1319ibus), .q(v1319obus), .dec(dec[1319]));
wire [data_w*2-1:0] v1320ibus;
wire [temp_w*2-1:0] v1320obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1320 (.l(l[1320*data_w +:data_w]), .r(v1320ibus), .q(v1320obus), .dec(dec[1320]));
wire [data_w*2-1:0] v1321ibus;
wire [temp_w*2-1:0] v1321obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1321 (.l(l[1321*data_w +:data_w]), .r(v1321ibus), .q(v1321obus), .dec(dec[1321]));
wire [data_w*2-1:0] v1322ibus;
wire [temp_w*2-1:0] v1322obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1322 (.l(l[1322*data_w +:data_w]), .r(v1322ibus), .q(v1322obus), .dec(dec[1322]));
wire [data_w*2-1:0] v1323ibus;
wire [temp_w*2-1:0] v1323obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1323 (.l(l[1323*data_w +:data_w]), .r(v1323ibus), .q(v1323obus), .dec(dec[1323]));
wire [data_w*2-1:0] v1324ibus;
wire [temp_w*2-1:0] v1324obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1324 (.l(l[1324*data_w +:data_w]), .r(v1324ibus), .q(v1324obus), .dec(dec[1324]));
wire [data_w*2-1:0] v1325ibus;
wire [temp_w*2-1:0] v1325obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1325 (.l(l[1325*data_w +:data_w]), .r(v1325ibus), .q(v1325obus), .dec(dec[1325]));
wire [data_w*2-1:0] v1326ibus;
wire [temp_w*2-1:0] v1326obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1326 (.l(l[1326*data_w +:data_w]), .r(v1326ibus), .q(v1326obus), .dec(dec[1326]));
wire [data_w*2-1:0] v1327ibus;
wire [temp_w*2-1:0] v1327obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1327 (.l(l[1327*data_w +:data_w]), .r(v1327ibus), .q(v1327obus), .dec(dec[1327]));
wire [data_w*2-1:0] v1328ibus;
wire [temp_w*2-1:0] v1328obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1328 (.l(l[1328*data_w +:data_w]), .r(v1328ibus), .q(v1328obus), .dec(dec[1328]));
wire [data_w*2-1:0] v1329ibus;
wire [temp_w*2-1:0] v1329obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1329 (.l(l[1329*data_w +:data_w]), .r(v1329ibus), .q(v1329obus), .dec(dec[1329]));
wire [data_w*2-1:0] v1330ibus;
wire [temp_w*2-1:0] v1330obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1330 (.l(l[1330*data_w +:data_w]), .r(v1330ibus), .q(v1330obus), .dec(dec[1330]));
wire [data_w*2-1:0] v1331ibus;
wire [temp_w*2-1:0] v1331obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1331 (.l(l[1331*data_w +:data_w]), .r(v1331ibus), .q(v1331obus), .dec(dec[1331]));
wire [data_w*2-1:0] v1332ibus;
wire [temp_w*2-1:0] v1332obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1332 (.l(l[1332*data_w +:data_w]), .r(v1332ibus), .q(v1332obus), .dec(dec[1332]));
wire [data_w*2-1:0] v1333ibus;
wire [temp_w*2-1:0] v1333obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1333 (.l(l[1333*data_w +:data_w]), .r(v1333ibus), .q(v1333obus), .dec(dec[1333]));
wire [data_w*2-1:0] v1334ibus;
wire [temp_w*2-1:0] v1334obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1334 (.l(l[1334*data_w +:data_w]), .r(v1334ibus), .q(v1334obus), .dec(dec[1334]));
wire [data_w*2-1:0] v1335ibus;
wire [temp_w*2-1:0] v1335obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1335 (.l(l[1335*data_w +:data_w]), .r(v1335ibus), .q(v1335obus), .dec(dec[1335]));
wire [data_w*2-1:0] v1336ibus;
wire [temp_w*2-1:0] v1336obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1336 (.l(l[1336*data_w +:data_w]), .r(v1336ibus), .q(v1336obus), .dec(dec[1336]));
wire [data_w*2-1:0] v1337ibus;
wire [temp_w*2-1:0] v1337obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1337 (.l(l[1337*data_w +:data_w]), .r(v1337ibus), .q(v1337obus), .dec(dec[1337]));
wire [data_w*2-1:0] v1338ibus;
wire [temp_w*2-1:0] v1338obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1338 (.l(l[1338*data_w +:data_w]), .r(v1338ibus), .q(v1338obus), .dec(dec[1338]));
wire [data_w*2-1:0] v1339ibus;
wire [temp_w*2-1:0] v1339obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1339 (.l(l[1339*data_w +:data_w]), .r(v1339ibus), .q(v1339obus), .dec(dec[1339]));
wire [data_w*2-1:0] v1340ibus;
wire [temp_w*2-1:0] v1340obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1340 (.l(l[1340*data_w +:data_w]), .r(v1340ibus), .q(v1340obus), .dec(dec[1340]));
wire [data_w*2-1:0] v1341ibus;
wire [temp_w*2-1:0] v1341obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1341 (.l(l[1341*data_w +:data_w]), .r(v1341ibus), .q(v1341obus), .dec(dec[1341]));
wire [data_w*2-1:0] v1342ibus;
wire [temp_w*2-1:0] v1342obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1342 (.l(l[1342*data_w +:data_w]), .r(v1342ibus), .q(v1342obus), .dec(dec[1342]));
wire [data_w*2-1:0] v1343ibus;
wire [temp_w*2-1:0] v1343obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1343 (.l(l[1343*data_w +:data_w]), .r(v1343ibus), .q(v1343obus), .dec(dec[1343]));
wire [data_w*2-1:0] v1344ibus;
wire [temp_w*2-1:0] v1344obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1344 (.l(l[1344*data_w +:data_w]), .r(v1344ibus), .q(v1344obus), .dec(dec[1344]));
wire [data_w*2-1:0] v1345ibus;
wire [temp_w*2-1:0] v1345obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1345 (.l(l[1345*data_w +:data_w]), .r(v1345ibus), .q(v1345obus), .dec(dec[1345]));
wire [data_w*2-1:0] v1346ibus;
wire [temp_w*2-1:0] v1346obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1346 (.l(l[1346*data_w +:data_w]), .r(v1346ibus), .q(v1346obus), .dec(dec[1346]));
wire [data_w*2-1:0] v1347ibus;
wire [temp_w*2-1:0] v1347obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1347 (.l(l[1347*data_w +:data_w]), .r(v1347ibus), .q(v1347obus), .dec(dec[1347]));
wire [data_w*2-1:0] v1348ibus;
wire [temp_w*2-1:0] v1348obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1348 (.l(l[1348*data_w +:data_w]), .r(v1348ibus), .q(v1348obus), .dec(dec[1348]));
wire [data_w*2-1:0] v1349ibus;
wire [temp_w*2-1:0] v1349obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1349 (.l(l[1349*data_w +:data_w]), .r(v1349ibus), .q(v1349obus), .dec(dec[1349]));
wire [data_w*2-1:0] v1350ibus;
wire [temp_w*2-1:0] v1350obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1350 (.l(l[1350*data_w +:data_w]), .r(v1350ibus), .q(v1350obus), .dec(dec[1350]));
wire [data_w*2-1:0] v1351ibus;
wire [temp_w*2-1:0] v1351obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1351 (.l(l[1351*data_w +:data_w]), .r(v1351ibus), .q(v1351obus), .dec(dec[1351]));
wire [data_w*2-1:0] v1352ibus;
wire [temp_w*2-1:0] v1352obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1352 (.l(l[1352*data_w +:data_w]), .r(v1352ibus), .q(v1352obus), .dec(dec[1352]));
wire [data_w*2-1:0] v1353ibus;
wire [temp_w*2-1:0] v1353obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1353 (.l(l[1353*data_w +:data_w]), .r(v1353ibus), .q(v1353obus), .dec(dec[1353]));
wire [data_w*2-1:0] v1354ibus;
wire [temp_w*2-1:0] v1354obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1354 (.l(l[1354*data_w +:data_w]), .r(v1354ibus), .q(v1354obus), .dec(dec[1354]));
wire [data_w*2-1:0] v1355ibus;
wire [temp_w*2-1:0] v1355obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1355 (.l(l[1355*data_w +:data_w]), .r(v1355ibus), .q(v1355obus), .dec(dec[1355]));
wire [data_w*2-1:0] v1356ibus;
wire [temp_w*2-1:0] v1356obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1356 (.l(l[1356*data_w +:data_w]), .r(v1356ibus), .q(v1356obus), .dec(dec[1356]));
wire [data_w*2-1:0] v1357ibus;
wire [temp_w*2-1:0] v1357obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1357 (.l(l[1357*data_w +:data_w]), .r(v1357ibus), .q(v1357obus), .dec(dec[1357]));
wire [data_w*2-1:0] v1358ibus;
wire [temp_w*2-1:0] v1358obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1358 (.l(l[1358*data_w +:data_w]), .r(v1358ibus), .q(v1358obus), .dec(dec[1358]));
wire [data_w*2-1:0] v1359ibus;
wire [temp_w*2-1:0] v1359obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1359 (.l(l[1359*data_w +:data_w]), .r(v1359ibus), .q(v1359obus), .dec(dec[1359]));
wire [data_w*2-1:0] v1360ibus;
wire [temp_w*2-1:0] v1360obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1360 (.l(l[1360*data_w +:data_w]), .r(v1360ibus), .q(v1360obus), .dec(dec[1360]));
wire [data_w*2-1:0] v1361ibus;
wire [temp_w*2-1:0] v1361obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1361 (.l(l[1361*data_w +:data_w]), .r(v1361ibus), .q(v1361obus), .dec(dec[1361]));
wire [data_w*2-1:0] v1362ibus;
wire [temp_w*2-1:0] v1362obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1362 (.l(l[1362*data_w +:data_w]), .r(v1362ibus), .q(v1362obus), .dec(dec[1362]));
wire [data_w*2-1:0] v1363ibus;
wire [temp_w*2-1:0] v1363obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1363 (.l(l[1363*data_w +:data_w]), .r(v1363ibus), .q(v1363obus), .dec(dec[1363]));
wire [data_w*2-1:0] v1364ibus;
wire [temp_w*2-1:0] v1364obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1364 (.l(l[1364*data_w +:data_w]), .r(v1364ibus), .q(v1364obus), .dec(dec[1364]));
wire [data_w*2-1:0] v1365ibus;
wire [temp_w*2-1:0] v1365obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1365 (.l(l[1365*data_w +:data_w]), .r(v1365ibus), .q(v1365obus), .dec(dec[1365]));
wire [data_w*2-1:0] v1366ibus;
wire [temp_w*2-1:0] v1366obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1366 (.l(l[1366*data_w +:data_w]), .r(v1366ibus), .q(v1366obus), .dec(dec[1366]));
wire [data_w*2-1:0] v1367ibus;
wire [temp_w*2-1:0] v1367obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1367 (.l(l[1367*data_w +:data_w]), .r(v1367ibus), .q(v1367obus), .dec(dec[1367]));
wire [data_w*2-1:0] v1368ibus;
wire [temp_w*2-1:0] v1368obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1368 (.l(l[1368*data_w +:data_w]), .r(v1368ibus), .q(v1368obus), .dec(dec[1368]));
wire [data_w*2-1:0] v1369ibus;
wire [temp_w*2-1:0] v1369obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1369 (.l(l[1369*data_w +:data_w]), .r(v1369ibus), .q(v1369obus), .dec(dec[1369]));
wire [data_w*2-1:0] v1370ibus;
wire [temp_w*2-1:0] v1370obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1370 (.l(l[1370*data_w +:data_w]), .r(v1370ibus), .q(v1370obus), .dec(dec[1370]));
wire [data_w*2-1:0] v1371ibus;
wire [temp_w*2-1:0] v1371obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1371 (.l(l[1371*data_w +:data_w]), .r(v1371ibus), .q(v1371obus), .dec(dec[1371]));
wire [data_w*2-1:0] v1372ibus;
wire [temp_w*2-1:0] v1372obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1372 (.l(l[1372*data_w +:data_w]), .r(v1372ibus), .q(v1372obus), .dec(dec[1372]));
wire [data_w*2-1:0] v1373ibus;
wire [temp_w*2-1:0] v1373obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1373 (.l(l[1373*data_w +:data_w]), .r(v1373ibus), .q(v1373obus), .dec(dec[1373]));
wire [data_w*2-1:0] v1374ibus;
wire [temp_w*2-1:0] v1374obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1374 (.l(l[1374*data_w +:data_w]), .r(v1374ibus), .q(v1374obus), .dec(dec[1374]));
wire [data_w*2-1:0] v1375ibus;
wire [temp_w*2-1:0] v1375obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1375 (.l(l[1375*data_w +:data_w]), .r(v1375ibus), .q(v1375obus), .dec(dec[1375]));
wire [data_w*2-1:0] v1376ibus;
wire [temp_w*2-1:0] v1376obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1376 (.l(l[1376*data_w +:data_w]), .r(v1376ibus), .q(v1376obus), .dec(dec[1376]));
wire [data_w*2-1:0] v1377ibus;
wire [temp_w*2-1:0] v1377obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1377 (.l(l[1377*data_w +:data_w]), .r(v1377ibus), .q(v1377obus), .dec(dec[1377]));
wire [data_w*2-1:0] v1378ibus;
wire [temp_w*2-1:0] v1378obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1378 (.l(l[1378*data_w +:data_w]), .r(v1378ibus), .q(v1378obus), .dec(dec[1378]));
wire [data_w*2-1:0] v1379ibus;
wire [temp_w*2-1:0] v1379obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1379 (.l(l[1379*data_w +:data_w]), .r(v1379ibus), .q(v1379obus), .dec(dec[1379]));
wire [data_w*2-1:0] v1380ibus;
wire [temp_w*2-1:0] v1380obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1380 (.l(l[1380*data_w +:data_w]), .r(v1380ibus), .q(v1380obus), .dec(dec[1380]));
wire [data_w*2-1:0] v1381ibus;
wire [temp_w*2-1:0] v1381obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1381 (.l(l[1381*data_w +:data_w]), .r(v1381ibus), .q(v1381obus), .dec(dec[1381]));
wire [data_w*2-1:0] v1382ibus;
wire [temp_w*2-1:0] v1382obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1382 (.l(l[1382*data_w +:data_w]), .r(v1382ibus), .q(v1382obus), .dec(dec[1382]));
wire [data_w*2-1:0] v1383ibus;
wire [temp_w*2-1:0] v1383obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1383 (.l(l[1383*data_w +:data_w]), .r(v1383ibus), .q(v1383obus), .dec(dec[1383]));
wire [data_w*2-1:0] v1384ibus;
wire [temp_w*2-1:0] v1384obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1384 (.l(l[1384*data_w +:data_w]), .r(v1384ibus), .q(v1384obus), .dec(dec[1384]));
wire [data_w*2-1:0] v1385ibus;
wire [temp_w*2-1:0] v1385obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1385 (.l(l[1385*data_w +:data_w]), .r(v1385ibus), .q(v1385obus), .dec(dec[1385]));
wire [data_w*2-1:0] v1386ibus;
wire [temp_w*2-1:0] v1386obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1386 (.l(l[1386*data_w +:data_w]), .r(v1386ibus), .q(v1386obus), .dec(dec[1386]));
wire [data_w*2-1:0] v1387ibus;
wire [temp_w*2-1:0] v1387obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1387 (.l(l[1387*data_w +:data_w]), .r(v1387ibus), .q(v1387obus), .dec(dec[1387]));
wire [data_w*2-1:0] v1388ibus;
wire [temp_w*2-1:0] v1388obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1388 (.l(l[1388*data_w +:data_w]), .r(v1388ibus), .q(v1388obus), .dec(dec[1388]));
wire [data_w*2-1:0] v1389ibus;
wire [temp_w*2-1:0] v1389obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1389 (.l(l[1389*data_w +:data_w]), .r(v1389ibus), .q(v1389obus), .dec(dec[1389]));
wire [data_w*2-1:0] v1390ibus;
wire [temp_w*2-1:0] v1390obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1390 (.l(l[1390*data_w +:data_w]), .r(v1390ibus), .q(v1390obus), .dec(dec[1390]));
wire [data_w*2-1:0] v1391ibus;
wire [temp_w*2-1:0] v1391obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1391 (.l(l[1391*data_w +:data_w]), .r(v1391ibus), .q(v1391obus), .dec(dec[1391]));
wire [data_w*2-1:0] v1392ibus;
wire [temp_w*2-1:0] v1392obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1392 (.l(l[1392*data_w +:data_w]), .r(v1392ibus), .q(v1392obus), .dec(dec[1392]));
wire [data_w*2-1:0] v1393ibus;
wire [temp_w*2-1:0] v1393obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1393 (.l(l[1393*data_w +:data_w]), .r(v1393ibus), .q(v1393obus), .dec(dec[1393]));
wire [data_w*2-1:0] v1394ibus;
wire [temp_w*2-1:0] v1394obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1394 (.l(l[1394*data_w +:data_w]), .r(v1394ibus), .q(v1394obus), .dec(dec[1394]));
wire [data_w*2-1:0] v1395ibus;
wire [temp_w*2-1:0] v1395obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1395 (.l(l[1395*data_w +:data_w]), .r(v1395ibus), .q(v1395obus), .dec(dec[1395]));
wire [data_w*2-1:0] v1396ibus;
wire [temp_w*2-1:0] v1396obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1396 (.l(l[1396*data_w +:data_w]), .r(v1396ibus), .q(v1396obus), .dec(dec[1396]));
wire [data_w*2-1:0] v1397ibus;
wire [temp_w*2-1:0] v1397obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1397 (.l(l[1397*data_w +:data_w]), .r(v1397ibus), .q(v1397obus), .dec(dec[1397]));
wire [data_w*2-1:0] v1398ibus;
wire [temp_w*2-1:0] v1398obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1398 (.l(l[1398*data_w +:data_w]), .r(v1398ibus), .q(v1398obus), .dec(dec[1398]));
wire [data_w*2-1:0] v1399ibus;
wire [temp_w*2-1:0] v1399obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1399 (.l(l[1399*data_w +:data_w]), .r(v1399ibus), .q(v1399obus), .dec(dec[1399]));
wire [data_w*2-1:0] v1400ibus;
wire [temp_w*2-1:0] v1400obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1400 (.l(l[1400*data_w +:data_w]), .r(v1400ibus), .q(v1400obus), .dec(dec[1400]));
wire [data_w*2-1:0] v1401ibus;
wire [temp_w*2-1:0] v1401obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1401 (.l(l[1401*data_w +:data_w]), .r(v1401ibus), .q(v1401obus), .dec(dec[1401]));
wire [data_w*2-1:0] v1402ibus;
wire [temp_w*2-1:0] v1402obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1402 (.l(l[1402*data_w +:data_w]), .r(v1402ibus), .q(v1402obus), .dec(dec[1402]));
wire [data_w*2-1:0] v1403ibus;
wire [temp_w*2-1:0] v1403obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1403 (.l(l[1403*data_w +:data_w]), .r(v1403ibus), .q(v1403obus), .dec(dec[1403]));
wire [data_w*2-1:0] v1404ibus;
wire [temp_w*2-1:0] v1404obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1404 (.l(l[1404*data_w +:data_w]), .r(v1404ibus), .q(v1404obus), .dec(dec[1404]));
wire [data_w*2-1:0] v1405ibus;
wire [temp_w*2-1:0] v1405obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1405 (.l(l[1405*data_w +:data_w]), .r(v1405ibus), .q(v1405obus), .dec(dec[1405]));
wire [data_w*2-1:0] v1406ibus;
wire [temp_w*2-1:0] v1406obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1406 (.l(l[1406*data_w +:data_w]), .r(v1406ibus), .q(v1406obus), .dec(dec[1406]));
wire [data_w*2-1:0] v1407ibus;
wire [temp_w*2-1:0] v1407obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1407 (.l(l[1407*data_w +:data_w]), .r(v1407ibus), .q(v1407obus), .dec(dec[1407]));
wire [data_w*2-1:0] v1408ibus;
wire [temp_w*2-1:0] v1408obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1408 (.l(l[1408*data_w +:data_w]), .r(v1408ibus), .q(v1408obus), .dec(dec[1408]));
wire [data_w*2-1:0] v1409ibus;
wire [temp_w*2-1:0] v1409obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1409 (.l(l[1409*data_w +:data_w]), .r(v1409ibus), .q(v1409obus), .dec(dec[1409]));
wire [data_w*2-1:0] v1410ibus;
wire [temp_w*2-1:0] v1410obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1410 (.l(l[1410*data_w +:data_w]), .r(v1410ibus), .q(v1410obus), .dec(dec[1410]));
wire [data_w*2-1:0] v1411ibus;
wire [temp_w*2-1:0] v1411obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1411 (.l(l[1411*data_w +:data_w]), .r(v1411ibus), .q(v1411obus), .dec(dec[1411]));
wire [data_w*2-1:0] v1412ibus;
wire [temp_w*2-1:0] v1412obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1412 (.l(l[1412*data_w +:data_w]), .r(v1412ibus), .q(v1412obus), .dec(dec[1412]));
wire [data_w*2-1:0] v1413ibus;
wire [temp_w*2-1:0] v1413obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1413 (.l(l[1413*data_w +:data_w]), .r(v1413ibus), .q(v1413obus), .dec(dec[1413]));
wire [data_w*2-1:0] v1414ibus;
wire [temp_w*2-1:0] v1414obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1414 (.l(l[1414*data_w +:data_w]), .r(v1414ibus), .q(v1414obus), .dec(dec[1414]));
wire [data_w*2-1:0] v1415ibus;
wire [temp_w*2-1:0] v1415obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1415 (.l(l[1415*data_w +:data_w]), .r(v1415ibus), .q(v1415obus), .dec(dec[1415]));
wire [data_w*2-1:0] v1416ibus;
wire [temp_w*2-1:0] v1416obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1416 (.l(l[1416*data_w +:data_w]), .r(v1416ibus), .q(v1416obus), .dec(dec[1416]));
wire [data_w*2-1:0] v1417ibus;
wire [temp_w*2-1:0] v1417obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1417 (.l(l[1417*data_w +:data_w]), .r(v1417ibus), .q(v1417obus), .dec(dec[1417]));
wire [data_w*2-1:0] v1418ibus;
wire [temp_w*2-1:0] v1418obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1418 (.l(l[1418*data_w +:data_w]), .r(v1418ibus), .q(v1418obus), .dec(dec[1418]));
wire [data_w*2-1:0] v1419ibus;
wire [temp_w*2-1:0] v1419obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1419 (.l(l[1419*data_w +:data_w]), .r(v1419ibus), .q(v1419obus), .dec(dec[1419]));
wire [data_w*2-1:0] v1420ibus;
wire [temp_w*2-1:0] v1420obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1420 (.l(l[1420*data_w +:data_w]), .r(v1420ibus), .q(v1420obus), .dec(dec[1420]));
wire [data_w*2-1:0] v1421ibus;
wire [temp_w*2-1:0] v1421obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1421 (.l(l[1421*data_w +:data_w]), .r(v1421ibus), .q(v1421obus), .dec(dec[1421]));
wire [data_w*2-1:0] v1422ibus;
wire [temp_w*2-1:0] v1422obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1422 (.l(l[1422*data_w +:data_w]), .r(v1422ibus), .q(v1422obus), .dec(dec[1422]));
wire [data_w*2-1:0] v1423ibus;
wire [temp_w*2-1:0] v1423obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1423 (.l(l[1423*data_w +:data_w]), .r(v1423ibus), .q(v1423obus), .dec(dec[1423]));
wire [data_w*2-1:0] v1424ibus;
wire [temp_w*2-1:0] v1424obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1424 (.l(l[1424*data_w +:data_w]), .r(v1424ibus), .q(v1424obus), .dec(dec[1424]));
wire [data_w*2-1:0] v1425ibus;
wire [temp_w*2-1:0] v1425obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1425 (.l(l[1425*data_w +:data_w]), .r(v1425ibus), .q(v1425obus), .dec(dec[1425]));
wire [data_w*2-1:0] v1426ibus;
wire [temp_w*2-1:0] v1426obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1426 (.l(l[1426*data_w +:data_w]), .r(v1426ibus), .q(v1426obus), .dec(dec[1426]));
wire [data_w*2-1:0] v1427ibus;
wire [temp_w*2-1:0] v1427obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1427 (.l(l[1427*data_w +:data_w]), .r(v1427ibus), .q(v1427obus), .dec(dec[1427]));
wire [data_w*2-1:0] v1428ibus;
wire [temp_w*2-1:0] v1428obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1428 (.l(l[1428*data_w +:data_w]), .r(v1428ibus), .q(v1428obus), .dec(dec[1428]));
wire [data_w*2-1:0] v1429ibus;
wire [temp_w*2-1:0] v1429obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1429 (.l(l[1429*data_w +:data_w]), .r(v1429ibus), .q(v1429obus), .dec(dec[1429]));
wire [data_w*2-1:0] v1430ibus;
wire [temp_w*2-1:0] v1430obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1430 (.l(l[1430*data_w +:data_w]), .r(v1430ibus), .q(v1430obus), .dec(dec[1430]));
wire [data_w*2-1:0] v1431ibus;
wire [temp_w*2-1:0] v1431obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1431 (.l(l[1431*data_w +:data_w]), .r(v1431ibus), .q(v1431obus), .dec(dec[1431]));
wire [data_w*2-1:0] v1432ibus;
wire [temp_w*2-1:0] v1432obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1432 (.l(l[1432*data_w +:data_w]), .r(v1432ibus), .q(v1432obus), .dec(dec[1432]));
wire [data_w*2-1:0] v1433ibus;
wire [temp_w*2-1:0] v1433obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1433 (.l(l[1433*data_w +:data_w]), .r(v1433ibus), .q(v1433obus), .dec(dec[1433]));
wire [data_w*2-1:0] v1434ibus;
wire [temp_w*2-1:0] v1434obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1434 (.l(l[1434*data_w +:data_w]), .r(v1434ibus), .q(v1434obus), .dec(dec[1434]));
wire [data_w*2-1:0] v1435ibus;
wire [temp_w*2-1:0] v1435obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1435 (.l(l[1435*data_w +:data_w]), .r(v1435ibus), .q(v1435obus), .dec(dec[1435]));
wire [data_w*2-1:0] v1436ibus;
wire [temp_w*2-1:0] v1436obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1436 (.l(l[1436*data_w +:data_w]), .r(v1436ibus), .q(v1436obus), .dec(dec[1436]));
wire [data_w*2-1:0] v1437ibus;
wire [temp_w*2-1:0] v1437obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1437 (.l(l[1437*data_w +:data_w]), .r(v1437ibus), .q(v1437obus), .dec(dec[1437]));
wire [data_w*2-1:0] v1438ibus;
wire [temp_w*2-1:0] v1438obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1438 (.l(l[1438*data_w +:data_w]), .r(v1438ibus), .q(v1438obus), .dec(dec[1438]));
wire [data_w*2-1:0] v1439ibus;
wire [temp_w*2-1:0] v1439obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1439 (.l(l[1439*data_w +:data_w]), .r(v1439ibus), .q(v1439obus), .dec(dec[1439]));
wire [data_w*2-1:0] v1440ibus;
wire [temp_w*2-1:0] v1440obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1440 (.l(l[1440*data_w +:data_w]), .r(v1440ibus), .q(v1440obus), .dec(dec[1440]));
wire [data_w*2-1:0] v1441ibus;
wire [temp_w*2-1:0] v1441obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1441 (.l(l[1441*data_w +:data_w]), .r(v1441ibus), .q(v1441obus), .dec(dec[1441]));
wire [data_w*2-1:0] v1442ibus;
wire [temp_w*2-1:0] v1442obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1442 (.l(l[1442*data_w +:data_w]), .r(v1442ibus), .q(v1442obus), .dec(dec[1442]));
wire [data_w*2-1:0] v1443ibus;
wire [temp_w*2-1:0] v1443obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1443 (.l(l[1443*data_w +:data_w]), .r(v1443ibus), .q(v1443obus), .dec(dec[1443]));
wire [data_w*2-1:0] v1444ibus;
wire [temp_w*2-1:0] v1444obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1444 (.l(l[1444*data_w +:data_w]), .r(v1444ibus), .q(v1444obus), .dec(dec[1444]));
wire [data_w*2-1:0] v1445ibus;
wire [temp_w*2-1:0] v1445obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1445 (.l(l[1445*data_w +:data_w]), .r(v1445ibus), .q(v1445obus), .dec(dec[1445]));
wire [data_w*2-1:0] v1446ibus;
wire [temp_w*2-1:0] v1446obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1446 (.l(l[1446*data_w +:data_w]), .r(v1446ibus), .q(v1446obus), .dec(dec[1446]));
wire [data_w*2-1:0] v1447ibus;
wire [temp_w*2-1:0] v1447obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1447 (.l(l[1447*data_w +:data_w]), .r(v1447ibus), .q(v1447obus), .dec(dec[1447]));
wire [data_w*2-1:0] v1448ibus;
wire [temp_w*2-1:0] v1448obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1448 (.l(l[1448*data_w +:data_w]), .r(v1448ibus), .q(v1448obus), .dec(dec[1448]));
wire [data_w*2-1:0] v1449ibus;
wire [temp_w*2-1:0] v1449obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1449 (.l(l[1449*data_w +:data_w]), .r(v1449ibus), .q(v1449obus), .dec(dec[1449]));
wire [data_w*2-1:0] v1450ibus;
wire [temp_w*2-1:0] v1450obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1450 (.l(l[1450*data_w +:data_w]), .r(v1450ibus), .q(v1450obus), .dec(dec[1450]));
wire [data_w*2-1:0] v1451ibus;
wire [temp_w*2-1:0] v1451obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1451 (.l(l[1451*data_w +:data_w]), .r(v1451ibus), .q(v1451obus), .dec(dec[1451]));
wire [data_w*2-1:0] v1452ibus;
wire [temp_w*2-1:0] v1452obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1452 (.l(l[1452*data_w +:data_w]), .r(v1452ibus), .q(v1452obus), .dec(dec[1452]));
wire [data_w*2-1:0] v1453ibus;
wire [temp_w*2-1:0] v1453obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1453 (.l(l[1453*data_w +:data_w]), .r(v1453ibus), .q(v1453obus), .dec(dec[1453]));
wire [data_w*2-1:0] v1454ibus;
wire [temp_w*2-1:0] v1454obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1454 (.l(l[1454*data_w +:data_w]), .r(v1454ibus), .q(v1454obus), .dec(dec[1454]));
wire [data_w*2-1:0] v1455ibus;
wire [temp_w*2-1:0] v1455obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1455 (.l(l[1455*data_w +:data_w]), .r(v1455ibus), .q(v1455obus), .dec(dec[1455]));
wire [data_w*2-1:0] v1456ibus;
wire [temp_w*2-1:0] v1456obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1456 (.l(l[1456*data_w +:data_w]), .r(v1456ibus), .q(v1456obus), .dec(dec[1456]));
wire [data_w*2-1:0] v1457ibus;
wire [temp_w*2-1:0] v1457obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1457 (.l(l[1457*data_w +:data_w]), .r(v1457ibus), .q(v1457obus), .dec(dec[1457]));
wire [data_w*2-1:0] v1458ibus;
wire [temp_w*2-1:0] v1458obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1458 (.l(l[1458*data_w +:data_w]), .r(v1458ibus), .q(v1458obus), .dec(dec[1458]));
wire [data_w*2-1:0] v1459ibus;
wire [temp_w*2-1:0] v1459obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1459 (.l(l[1459*data_w +:data_w]), .r(v1459ibus), .q(v1459obus), .dec(dec[1459]));
wire [data_w*2-1:0] v1460ibus;
wire [temp_w*2-1:0] v1460obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1460 (.l(l[1460*data_w +:data_w]), .r(v1460ibus), .q(v1460obus), .dec(dec[1460]));
wire [data_w*2-1:0] v1461ibus;
wire [temp_w*2-1:0] v1461obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1461 (.l(l[1461*data_w +:data_w]), .r(v1461ibus), .q(v1461obus), .dec(dec[1461]));
wire [data_w*2-1:0] v1462ibus;
wire [temp_w*2-1:0] v1462obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1462 (.l(l[1462*data_w +:data_w]), .r(v1462ibus), .q(v1462obus), .dec(dec[1462]));
wire [data_w*2-1:0] v1463ibus;
wire [temp_w*2-1:0] v1463obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1463 (.l(l[1463*data_w +:data_w]), .r(v1463ibus), .q(v1463obus), .dec(dec[1463]));
wire [data_w*2-1:0] v1464ibus;
wire [temp_w*2-1:0] v1464obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1464 (.l(l[1464*data_w +:data_w]), .r(v1464ibus), .q(v1464obus), .dec(dec[1464]));
wire [data_w*2-1:0] v1465ibus;
wire [temp_w*2-1:0] v1465obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1465 (.l(l[1465*data_w +:data_w]), .r(v1465ibus), .q(v1465obus), .dec(dec[1465]));
wire [data_w*2-1:0] v1466ibus;
wire [temp_w*2-1:0] v1466obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1466 (.l(l[1466*data_w +:data_w]), .r(v1466ibus), .q(v1466obus), .dec(dec[1466]));
wire [data_w*2-1:0] v1467ibus;
wire [temp_w*2-1:0] v1467obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1467 (.l(l[1467*data_w +:data_w]), .r(v1467ibus), .q(v1467obus), .dec(dec[1467]));
wire [data_w*2-1:0] v1468ibus;
wire [temp_w*2-1:0] v1468obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1468 (.l(l[1468*data_w +:data_w]), .r(v1468ibus), .q(v1468obus), .dec(dec[1468]));
wire [data_w*2-1:0] v1469ibus;
wire [temp_w*2-1:0] v1469obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1469 (.l(l[1469*data_w +:data_w]), .r(v1469ibus), .q(v1469obus), .dec(dec[1469]));
wire [data_w*2-1:0] v1470ibus;
wire [temp_w*2-1:0] v1470obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1470 (.l(l[1470*data_w +:data_w]), .r(v1470ibus), .q(v1470obus), .dec(dec[1470]));
wire [data_w*2-1:0] v1471ibus;
wire [temp_w*2-1:0] v1471obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1471 (.l(l[1471*data_w +:data_w]), .r(v1471ibus), .q(v1471obus), .dec(dec[1471]));
wire [data_w*2-1:0] v1472ibus;
wire [temp_w*2-1:0] v1472obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1472 (.l(l[1472*data_w +:data_w]), .r(v1472ibus), .q(v1472obus), .dec(dec[1472]));
wire [data_w*2-1:0] v1473ibus;
wire [temp_w*2-1:0] v1473obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1473 (.l(l[1473*data_w +:data_w]), .r(v1473ibus), .q(v1473obus), .dec(dec[1473]));
wire [data_w*2-1:0] v1474ibus;
wire [temp_w*2-1:0] v1474obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1474 (.l(l[1474*data_w +:data_w]), .r(v1474ibus), .q(v1474obus), .dec(dec[1474]));
wire [data_w*2-1:0] v1475ibus;
wire [temp_w*2-1:0] v1475obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1475 (.l(l[1475*data_w +:data_w]), .r(v1475ibus), .q(v1475obus), .dec(dec[1475]));
wire [data_w*2-1:0] v1476ibus;
wire [temp_w*2-1:0] v1476obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1476 (.l(l[1476*data_w +:data_w]), .r(v1476ibus), .q(v1476obus), .dec(dec[1476]));
wire [data_w*2-1:0] v1477ibus;
wire [temp_w*2-1:0] v1477obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1477 (.l(l[1477*data_w +:data_w]), .r(v1477ibus), .q(v1477obus), .dec(dec[1477]));
wire [data_w*2-1:0] v1478ibus;
wire [temp_w*2-1:0] v1478obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1478 (.l(l[1478*data_w +:data_w]), .r(v1478ibus), .q(v1478obus), .dec(dec[1478]));
wire [data_w*2-1:0] v1479ibus;
wire [temp_w*2-1:0] v1479obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1479 (.l(l[1479*data_w +:data_w]), .r(v1479ibus), .q(v1479obus), .dec(dec[1479]));
wire [data_w*2-1:0] v1480ibus;
wire [temp_w*2-1:0] v1480obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1480 (.l(l[1480*data_w +:data_w]), .r(v1480ibus), .q(v1480obus), .dec(dec[1480]));
wire [data_w*2-1:0] v1481ibus;
wire [temp_w*2-1:0] v1481obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1481 (.l(l[1481*data_w +:data_w]), .r(v1481ibus), .q(v1481obus), .dec(dec[1481]));
wire [data_w*2-1:0] v1482ibus;
wire [temp_w*2-1:0] v1482obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1482 (.l(l[1482*data_w +:data_w]), .r(v1482ibus), .q(v1482obus), .dec(dec[1482]));
wire [data_w*2-1:0] v1483ibus;
wire [temp_w*2-1:0] v1483obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1483 (.l(l[1483*data_w +:data_w]), .r(v1483ibus), .q(v1483obus), .dec(dec[1483]));
wire [data_w*2-1:0] v1484ibus;
wire [temp_w*2-1:0] v1484obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1484 (.l(l[1484*data_w +:data_w]), .r(v1484ibus), .q(v1484obus), .dec(dec[1484]));
wire [data_w*2-1:0] v1485ibus;
wire [temp_w*2-1:0] v1485obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1485 (.l(l[1485*data_w +:data_w]), .r(v1485ibus), .q(v1485obus), .dec(dec[1485]));
wire [data_w*2-1:0] v1486ibus;
wire [temp_w*2-1:0] v1486obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1486 (.l(l[1486*data_w +:data_w]), .r(v1486ibus), .q(v1486obus), .dec(dec[1486]));
wire [data_w*2-1:0] v1487ibus;
wire [temp_w*2-1:0] v1487obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1487 (.l(l[1487*data_w +:data_w]), .r(v1487ibus), .q(v1487obus), .dec(dec[1487]));
wire [data_w*2-1:0] v1488ibus;
wire [temp_w*2-1:0] v1488obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1488 (.l(l[1488*data_w +:data_w]), .r(v1488ibus), .q(v1488obus), .dec(dec[1488]));
wire [data_w*2-1:0] v1489ibus;
wire [temp_w*2-1:0] v1489obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1489 (.l(l[1489*data_w +:data_w]), .r(v1489ibus), .q(v1489obus), .dec(dec[1489]));
wire [data_w*2-1:0] v1490ibus;
wire [temp_w*2-1:0] v1490obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1490 (.l(l[1490*data_w +:data_w]), .r(v1490ibus), .q(v1490obus), .dec(dec[1490]));
wire [data_w*2-1:0] v1491ibus;
wire [temp_w*2-1:0] v1491obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1491 (.l(l[1491*data_w +:data_w]), .r(v1491ibus), .q(v1491obus), .dec(dec[1491]));
wire [data_w*2-1:0] v1492ibus;
wire [temp_w*2-1:0] v1492obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1492 (.l(l[1492*data_w +:data_w]), .r(v1492ibus), .q(v1492obus), .dec(dec[1492]));
wire [data_w*2-1:0] v1493ibus;
wire [temp_w*2-1:0] v1493obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1493 (.l(l[1493*data_w +:data_w]), .r(v1493ibus), .q(v1493obus), .dec(dec[1493]));
wire [data_w*2-1:0] v1494ibus;
wire [temp_w*2-1:0] v1494obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1494 (.l(l[1494*data_w +:data_w]), .r(v1494ibus), .q(v1494obus), .dec(dec[1494]));
wire [data_w*2-1:0] v1495ibus;
wire [temp_w*2-1:0] v1495obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1495 (.l(l[1495*data_w +:data_w]), .r(v1495ibus), .q(v1495obus), .dec(dec[1495]));
wire [data_w*2-1:0] v1496ibus;
wire [temp_w*2-1:0] v1496obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1496 (.l(l[1496*data_w +:data_w]), .r(v1496ibus), .q(v1496obus), .dec(dec[1496]));
wire [data_w*2-1:0] v1497ibus;
wire [temp_w*2-1:0] v1497obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1497 (.l(l[1497*data_w +:data_w]), .r(v1497ibus), .q(v1497obus), .dec(dec[1497]));
wire [data_w*2-1:0] v1498ibus;
wire [temp_w*2-1:0] v1498obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1498 (.l(l[1498*data_w +:data_w]), .r(v1498ibus), .q(v1498obus), .dec(dec[1498]));
wire [data_w*2-1:0] v1499ibus;
wire [temp_w*2-1:0] v1499obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1499 (.l(l[1499*data_w +:data_w]), .r(v1499ibus), .q(v1499obus), .dec(dec[1499]));
wire [data_w*2-1:0] v1500ibus;
wire [temp_w*2-1:0] v1500obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1500 (.l(l[1500*data_w +:data_w]), .r(v1500ibus), .q(v1500obus), .dec(dec[1500]));
wire [data_w*2-1:0] v1501ibus;
wire [temp_w*2-1:0] v1501obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1501 (.l(l[1501*data_w +:data_w]), .r(v1501ibus), .q(v1501obus), .dec(dec[1501]));
wire [data_w*2-1:0] v1502ibus;
wire [temp_w*2-1:0] v1502obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1502 (.l(l[1502*data_w +:data_w]), .r(v1502ibus), .q(v1502obus), .dec(dec[1502]));
wire [data_w*2-1:0] v1503ibus;
wire [temp_w*2-1:0] v1503obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1503 (.l(l[1503*data_w +:data_w]), .r(v1503ibus), .q(v1503obus), .dec(dec[1503]));
wire [data_w*2-1:0] v1504ibus;
wire [temp_w*2-1:0] v1504obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1504 (.l(l[1504*data_w +:data_w]), .r(v1504ibus), .q(v1504obus), .dec(dec[1504]));
wire [data_w*2-1:0] v1505ibus;
wire [temp_w*2-1:0] v1505obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1505 (.l(l[1505*data_w +:data_w]), .r(v1505ibus), .q(v1505obus), .dec(dec[1505]));
wire [data_w*2-1:0] v1506ibus;
wire [temp_w*2-1:0] v1506obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1506 (.l(l[1506*data_w +:data_w]), .r(v1506ibus), .q(v1506obus), .dec(dec[1506]));
wire [data_w*2-1:0] v1507ibus;
wire [temp_w*2-1:0] v1507obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1507 (.l(l[1507*data_w +:data_w]), .r(v1507ibus), .q(v1507obus), .dec(dec[1507]));
wire [data_w*2-1:0] v1508ibus;
wire [temp_w*2-1:0] v1508obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1508 (.l(l[1508*data_w +:data_w]), .r(v1508ibus), .q(v1508obus), .dec(dec[1508]));
wire [data_w*2-1:0] v1509ibus;
wire [temp_w*2-1:0] v1509obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1509 (.l(l[1509*data_w +:data_w]), .r(v1509ibus), .q(v1509obus), .dec(dec[1509]));
wire [data_w*2-1:0] v1510ibus;
wire [temp_w*2-1:0] v1510obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1510 (.l(l[1510*data_w +:data_w]), .r(v1510ibus), .q(v1510obus), .dec(dec[1510]));
wire [data_w*2-1:0] v1511ibus;
wire [temp_w*2-1:0] v1511obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1511 (.l(l[1511*data_w +:data_w]), .r(v1511ibus), .q(v1511obus), .dec(dec[1511]));
wire [data_w*2-1:0] v1512ibus;
wire [temp_w*2-1:0] v1512obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1512 (.l(l[1512*data_w +:data_w]), .r(v1512ibus), .q(v1512obus), .dec(dec[1512]));
wire [data_w*2-1:0] v1513ibus;
wire [temp_w*2-1:0] v1513obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1513 (.l(l[1513*data_w +:data_w]), .r(v1513ibus), .q(v1513obus), .dec(dec[1513]));
wire [data_w*2-1:0] v1514ibus;
wire [temp_w*2-1:0] v1514obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1514 (.l(l[1514*data_w +:data_w]), .r(v1514ibus), .q(v1514obus), .dec(dec[1514]));
wire [data_w*2-1:0] v1515ibus;
wire [temp_w*2-1:0] v1515obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1515 (.l(l[1515*data_w +:data_w]), .r(v1515ibus), .q(v1515obus), .dec(dec[1515]));
wire [data_w*2-1:0] v1516ibus;
wire [temp_w*2-1:0] v1516obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1516 (.l(l[1516*data_w +:data_w]), .r(v1516ibus), .q(v1516obus), .dec(dec[1516]));
wire [data_w*2-1:0] v1517ibus;
wire [temp_w*2-1:0] v1517obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1517 (.l(l[1517*data_w +:data_w]), .r(v1517ibus), .q(v1517obus), .dec(dec[1517]));
wire [data_w*2-1:0] v1518ibus;
wire [temp_w*2-1:0] v1518obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1518 (.l(l[1518*data_w +:data_w]), .r(v1518ibus), .q(v1518obus), .dec(dec[1518]));
wire [data_w*2-1:0] v1519ibus;
wire [temp_w*2-1:0] v1519obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1519 (.l(l[1519*data_w +:data_w]), .r(v1519ibus), .q(v1519obus), .dec(dec[1519]));
wire [data_w*2-1:0] v1520ibus;
wire [temp_w*2-1:0] v1520obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1520 (.l(l[1520*data_w +:data_w]), .r(v1520ibus), .q(v1520obus), .dec(dec[1520]));
wire [data_w*2-1:0] v1521ibus;
wire [temp_w*2-1:0] v1521obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1521 (.l(l[1521*data_w +:data_w]), .r(v1521ibus), .q(v1521obus), .dec(dec[1521]));
wire [data_w*2-1:0] v1522ibus;
wire [temp_w*2-1:0] v1522obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1522 (.l(l[1522*data_w +:data_w]), .r(v1522ibus), .q(v1522obus), .dec(dec[1522]));
wire [data_w*2-1:0] v1523ibus;
wire [temp_w*2-1:0] v1523obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1523 (.l(l[1523*data_w +:data_w]), .r(v1523ibus), .q(v1523obus), .dec(dec[1523]));
wire [data_w*2-1:0] v1524ibus;
wire [temp_w*2-1:0] v1524obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1524 (.l(l[1524*data_w +:data_w]), .r(v1524ibus), .q(v1524obus), .dec(dec[1524]));
wire [data_w*2-1:0] v1525ibus;
wire [temp_w*2-1:0] v1525obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1525 (.l(l[1525*data_w +:data_w]), .r(v1525ibus), .q(v1525obus), .dec(dec[1525]));
wire [data_w*2-1:0] v1526ibus;
wire [temp_w*2-1:0] v1526obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1526 (.l(l[1526*data_w +:data_w]), .r(v1526ibus), .q(v1526obus), .dec(dec[1526]));
wire [data_w*2-1:0] v1527ibus;
wire [temp_w*2-1:0] v1527obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1527 (.l(l[1527*data_w +:data_w]), .r(v1527ibus), .q(v1527obus), .dec(dec[1527]));
wire [data_w*2-1:0] v1528ibus;
wire [temp_w*2-1:0] v1528obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1528 (.l(l[1528*data_w +:data_w]), .r(v1528ibus), .q(v1528obus), .dec(dec[1528]));
wire [data_w*2-1:0] v1529ibus;
wire [temp_w*2-1:0] v1529obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1529 (.l(l[1529*data_w +:data_w]), .r(v1529ibus), .q(v1529obus), .dec(dec[1529]));
wire [data_w*2-1:0] v1530ibus;
wire [temp_w*2-1:0] v1530obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1530 (.l(l[1530*data_w +:data_w]), .r(v1530ibus), .q(v1530obus), .dec(dec[1530]));
wire [data_w*2-1:0] v1531ibus;
wire [temp_w*2-1:0] v1531obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1531 (.l(l[1531*data_w +:data_w]), .r(v1531ibus), .q(v1531obus), .dec(dec[1531]));
wire [data_w*2-1:0] v1532ibus;
wire [temp_w*2-1:0] v1532obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1532 (.l(l[1532*data_w +:data_w]), .r(v1532ibus), .q(v1532obus), .dec(dec[1532]));
wire [data_w*2-1:0] v1533ibus;
wire [temp_w*2-1:0] v1533obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1533 (.l(l[1533*data_w +:data_w]), .r(v1533ibus), .q(v1533obus), .dec(dec[1533]));
wire [data_w*2-1:0] v1534ibus;
wire [temp_w*2-1:0] v1534obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1534 (.l(l[1534*data_w +:data_w]), .r(v1534ibus), .q(v1534obus), .dec(dec[1534]));
wire [data_w*2-1:0] v1535ibus;
wire [temp_w*2-1:0] v1535obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1535 (.l(l[1535*data_w +:data_w]), .r(v1535ibus), .q(v1535obus), .dec(dec[1535]));
wire [data_w*2-1:0] v1536ibus;
wire [temp_w*2-1:0] v1536obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1536 (.l(l[1536*data_w +:data_w]), .r(v1536ibus), .q(v1536obus), .dec(dec[1536]));
wire [data_w*2-1:0] v1537ibus;
wire [temp_w*2-1:0] v1537obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1537 (.l(l[1537*data_w +:data_w]), .r(v1537ibus), .q(v1537obus), .dec(dec[1537]));
wire [data_w*2-1:0] v1538ibus;
wire [temp_w*2-1:0] v1538obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1538 (.l(l[1538*data_w +:data_w]), .r(v1538ibus), .q(v1538obus), .dec(dec[1538]));
wire [data_w*2-1:0] v1539ibus;
wire [temp_w*2-1:0] v1539obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1539 (.l(l[1539*data_w +:data_w]), .r(v1539ibus), .q(v1539obus), .dec(dec[1539]));
wire [data_w*2-1:0] v1540ibus;
wire [temp_w*2-1:0] v1540obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1540 (.l(l[1540*data_w +:data_w]), .r(v1540ibus), .q(v1540obus), .dec(dec[1540]));
wire [data_w*2-1:0] v1541ibus;
wire [temp_w*2-1:0] v1541obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1541 (.l(l[1541*data_w +:data_w]), .r(v1541ibus), .q(v1541obus), .dec(dec[1541]));
wire [data_w*2-1:0] v1542ibus;
wire [temp_w*2-1:0] v1542obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1542 (.l(l[1542*data_w +:data_w]), .r(v1542ibus), .q(v1542obus), .dec(dec[1542]));
wire [data_w*2-1:0] v1543ibus;
wire [temp_w*2-1:0] v1543obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1543 (.l(l[1543*data_w +:data_w]), .r(v1543ibus), .q(v1543obus), .dec(dec[1543]));
wire [data_w*2-1:0] v1544ibus;
wire [temp_w*2-1:0] v1544obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1544 (.l(l[1544*data_w +:data_w]), .r(v1544ibus), .q(v1544obus), .dec(dec[1544]));
wire [data_w*2-1:0] v1545ibus;
wire [temp_w*2-1:0] v1545obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1545 (.l(l[1545*data_w +:data_w]), .r(v1545ibus), .q(v1545obus), .dec(dec[1545]));
wire [data_w*2-1:0] v1546ibus;
wire [temp_w*2-1:0] v1546obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1546 (.l(l[1546*data_w +:data_w]), .r(v1546ibus), .q(v1546obus), .dec(dec[1546]));
wire [data_w*2-1:0] v1547ibus;
wire [temp_w*2-1:0] v1547obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1547 (.l(l[1547*data_w +:data_w]), .r(v1547ibus), .q(v1547obus), .dec(dec[1547]));
wire [data_w*2-1:0] v1548ibus;
wire [temp_w*2-1:0] v1548obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1548 (.l(l[1548*data_w +:data_w]), .r(v1548ibus), .q(v1548obus), .dec(dec[1548]));
wire [data_w*2-1:0] v1549ibus;
wire [temp_w*2-1:0] v1549obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1549 (.l(l[1549*data_w +:data_w]), .r(v1549ibus), .q(v1549obus), .dec(dec[1549]));
wire [data_w*2-1:0] v1550ibus;
wire [temp_w*2-1:0] v1550obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1550 (.l(l[1550*data_w +:data_w]), .r(v1550ibus), .q(v1550obus), .dec(dec[1550]));
wire [data_w*2-1:0] v1551ibus;
wire [temp_w*2-1:0] v1551obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1551 (.l(l[1551*data_w +:data_w]), .r(v1551ibus), .q(v1551obus), .dec(dec[1551]));
wire [data_w*2-1:0] v1552ibus;
wire [temp_w*2-1:0] v1552obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1552 (.l(l[1552*data_w +:data_w]), .r(v1552ibus), .q(v1552obus), .dec(dec[1552]));
wire [data_w*2-1:0] v1553ibus;
wire [temp_w*2-1:0] v1553obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1553 (.l(l[1553*data_w +:data_w]), .r(v1553ibus), .q(v1553obus), .dec(dec[1553]));
wire [data_w*2-1:0] v1554ibus;
wire [temp_w*2-1:0] v1554obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1554 (.l(l[1554*data_w +:data_w]), .r(v1554ibus), .q(v1554obus), .dec(dec[1554]));
wire [data_w*2-1:0] v1555ibus;
wire [temp_w*2-1:0] v1555obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1555 (.l(l[1555*data_w +:data_w]), .r(v1555ibus), .q(v1555obus), .dec(dec[1555]));
wire [data_w*2-1:0] v1556ibus;
wire [temp_w*2-1:0] v1556obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1556 (.l(l[1556*data_w +:data_w]), .r(v1556ibus), .q(v1556obus), .dec(dec[1556]));
wire [data_w*2-1:0] v1557ibus;
wire [temp_w*2-1:0] v1557obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1557 (.l(l[1557*data_w +:data_w]), .r(v1557ibus), .q(v1557obus), .dec(dec[1557]));
wire [data_w*2-1:0] v1558ibus;
wire [temp_w*2-1:0] v1558obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1558 (.l(l[1558*data_w +:data_w]), .r(v1558ibus), .q(v1558obus), .dec(dec[1558]));
wire [data_w*2-1:0] v1559ibus;
wire [temp_w*2-1:0] v1559obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1559 (.l(l[1559*data_w +:data_w]), .r(v1559ibus), .q(v1559obus), .dec(dec[1559]));
wire [data_w*2-1:0] v1560ibus;
wire [temp_w*2-1:0] v1560obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1560 (.l(l[1560*data_w +:data_w]), .r(v1560ibus), .q(v1560obus), .dec(dec[1560]));
wire [data_w*2-1:0] v1561ibus;
wire [temp_w*2-1:0] v1561obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1561 (.l(l[1561*data_w +:data_w]), .r(v1561ibus), .q(v1561obus), .dec(dec[1561]));
wire [data_w*2-1:0] v1562ibus;
wire [temp_w*2-1:0] v1562obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1562 (.l(l[1562*data_w +:data_w]), .r(v1562ibus), .q(v1562obus), .dec(dec[1562]));
wire [data_w*2-1:0] v1563ibus;
wire [temp_w*2-1:0] v1563obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1563 (.l(l[1563*data_w +:data_w]), .r(v1563ibus), .q(v1563obus), .dec(dec[1563]));
wire [data_w*2-1:0] v1564ibus;
wire [temp_w*2-1:0] v1564obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1564 (.l(l[1564*data_w +:data_w]), .r(v1564ibus), .q(v1564obus), .dec(dec[1564]));
wire [data_w*2-1:0] v1565ibus;
wire [temp_w*2-1:0] v1565obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1565 (.l(l[1565*data_w +:data_w]), .r(v1565ibus), .q(v1565obus), .dec(dec[1565]));
wire [data_w*2-1:0] v1566ibus;
wire [temp_w*2-1:0] v1566obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1566 (.l(l[1566*data_w +:data_w]), .r(v1566ibus), .q(v1566obus), .dec(dec[1566]));
wire [data_w*2-1:0] v1567ibus;
wire [temp_w*2-1:0] v1567obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1567 (.l(l[1567*data_w +:data_w]), .r(v1567ibus), .q(v1567obus), .dec(dec[1567]));
wire [data_w*2-1:0] v1568ibus;
wire [temp_w*2-1:0] v1568obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1568 (.l(l[1568*data_w +:data_w]), .r(v1568ibus), .q(v1568obus), .dec(dec[1568]));
wire [data_w*2-1:0] v1569ibus;
wire [temp_w*2-1:0] v1569obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1569 (.l(l[1569*data_w +:data_w]), .r(v1569ibus), .q(v1569obus), .dec(dec[1569]));
wire [data_w*2-1:0] v1570ibus;
wire [temp_w*2-1:0] v1570obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1570 (.l(l[1570*data_w +:data_w]), .r(v1570ibus), .q(v1570obus), .dec(dec[1570]));
wire [data_w*2-1:0] v1571ibus;
wire [temp_w*2-1:0] v1571obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1571 (.l(l[1571*data_w +:data_w]), .r(v1571ibus), .q(v1571obus), .dec(dec[1571]));
wire [data_w*2-1:0] v1572ibus;
wire [temp_w*2-1:0] v1572obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1572 (.l(l[1572*data_w +:data_w]), .r(v1572ibus), .q(v1572obus), .dec(dec[1572]));
wire [data_w*2-1:0] v1573ibus;
wire [temp_w*2-1:0] v1573obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1573 (.l(l[1573*data_w +:data_w]), .r(v1573ibus), .q(v1573obus), .dec(dec[1573]));
wire [data_w*2-1:0] v1574ibus;
wire [temp_w*2-1:0] v1574obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1574 (.l(l[1574*data_w +:data_w]), .r(v1574ibus), .q(v1574obus), .dec(dec[1574]));
wire [data_w*2-1:0] v1575ibus;
wire [temp_w*2-1:0] v1575obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1575 (.l(l[1575*data_w +:data_w]), .r(v1575ibus), .q(v1575obus), .dec(dec[1575]));
wire [data_w*2-1:0] v1576ibus;
wire [temp_w*2-1:0] v1576obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1576 (.l(l[1576*data_w +:data_w]), .r(v1576ibus), .q(v1576obus), .dec(dec[1576]));
wire [data_w*2-1:0] v1577ibus;
wire [temp_w*2-1:0] v1577obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1577 (.l(l[1577*data_w +:data_w]), .r(v1577ibus), .q(v1577obus), .dec(dec[1577]));
wire [data_w*2-1:0] v1578ibus;
wire [temp_w*2-1:0] v1578obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1578 (.l(l[1578*data_w +:data_w]), .r(v1578ibus), .q(v1578obus), .dec(dec[1578]));
wire [data_w*2-1:0] v1579ibus;
wire [temp_w*2-1:0] v1579obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1579 (.l(l[1579*data_w +:data_w]), .r(v1579ibus), .q(v1579obus), .dec(dec[1579]));
wire [data_w*2-1:0] v1580ibus;
wire [temp_w*2-1:0] v1580obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1580 (.l(l[1580*data_w +:data_w]), .r(v1580ibus), .q(v1580obus), .dec(dec[1580]));
wire [data_w*2-1:0] v1581ibus;
wire [temp_w*2-1:0] v1581obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1581 (.l(l[1581*data_w +:data_w]), .r(v1581ibus), .q(v1581obus), .dec(dec[1581]));
wire [data_w*2-1:0] v1582ibus;
wire [temp_w*2-1:0] v1582obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1582 (.l(l[1582*data_w +:data_w]), .r(v1582ibus), .q(v1582obus), .dec(dec[1582]));
wire [data_w*2-1:0] v1583ibus;
wire [temp_w*2-1:0] v1583obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1583 (.l(l[1583*data_w +:data_w]), .r(v1583ibus), .q(v1583obus), .dec(dec[1583]));
wire [data_w*2-1:0] v1584ibus;
wire [temp_w*2-1:0] v1584obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1584 (.l(l[1584*data_w +:data_w]), .r(v1584ibus), .q(v1584obus), .dec(dec[1584]));
wire [data_w*2-1:0] v1585ibus;
wire [temp_w*2-1:0] v1585obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1585 (.l(l[1585*data_w +:data_w]), .r(v1585ibus), .q(v1585obus), .dec(dec[1585]));
wire [data_w*2-1:0] v1586ibus;
wire [temp_w*2-1:0] v1586obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1586 (.l(l[1586*data_w +:data_w]), .r(v1586ibus), .q(v1586obus), .dec(dec[1586]));
wire [data_w*2-1:0] v1587ibus;
wire [temp_w*2-1:0] v1587obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1587 (.l(l[1587*data_w +:data_w]), .r(v1587ibus), .q(v1587obus), .dec(dec[1587]));
wire [data_w*2-1:0] v1588ibus;
wire [temp_w*2-1:0] v1588obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1588 (.l(l[1588*data_w +:data_w]), .r(v1588ibus), .q(v1588obus), .dec(dec[1588]));
wire [data_w*2-1:0] v1589ibus;
wire [temp_w*2-1:0] v1589obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1589 (.l(l[1589*data_w +:data_w]), .r(v1589ibus), .q(v1589obus), .dec(dec[1589]));
wire [data_w*2-1:0] v1590ibus;
wire [temp_w*2-1:0] v1590obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1590 (.l(l[1590*data_w +:data_w]), .r(v1590ibus), .q(v1590obus), .dec(dec[1590]));
wire [data_w*2-1:0] v1591ibus;
wire [temp_w*2-1:0] v1591obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1591 (.l(l[1591*data_w +:data_w]), .r(v1591ibus), .q(v1591obus), .dec(dec[1591]));
wire [data_w*2-1:0] v1592ibus;
wire [temp_w*2-1:0] v1592obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1592 (.l(l[1592*data_w +:data_w]), .r(v1592ibus), .q(v1592obus), .dec(dec[1592]));
wire [data_w*2-1:0] v1593ibus;
wire [temp_w*2-1:0] v1593obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1593 (.l(l[1593*data_w +:data_w]), .r(v1593ibus), .q(v1593obus), .dec(dec[1593]));
wire [data_w*2-1:0] v1594ibus;
wire [temp_w*2-1:0] v1594obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1594 (.l(l[1594*data_w +:data_w]), .r(v1594ibus), .q(v1594obus), .dec(dec[1594]));
wire [data_w*2-1:0] v1595ibus;
wire [temp_w*2-1:0] v1595obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1595 (.l(l[1595*data_w +:data_w]), .r(v1595ibus), .q(v1595obus), .dec(dec[1595]));
wire [data_w*2-1:0] v1596ibus;
wire [temp_w*2-1:0] v1596obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1596 (.l(l[1596*data_w +:data_w]), .r(v1596ibus), .q(v1596obus), .dec(dec[1596]));
wire [data_w*2-1:0] v1597ibus;
wire [temp_w*2-1:0] v1597obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1597 (.l(l[1597*data_w +:data_w]), .r(v1597ibus), .q(v1597obus), .dec(dec[1597]));
wire [data_w*2-1:0] v1598ibus;
wire [temp_w*2-1:0] v1598obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1598 (.l(l[1598*data_w +:data_w]), .r(v1598ibus), .q(v1598obus), .dec(dec[1598]));
wire [data_w*2-1:0] v1599ibus;
wire [temp_w*2-1:0] v1599obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1599 (.l(l[1599*data_w +:data_w]), .r(v1599ibus), .q(v1599obus), .dec(dec[1599]));
wire [data_w*2-1:0] v1600ibus;
wire [temp_w*2-1:0] v1600obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1600 (.l(l[1600*data_w +:data_w]), .r(v1600ibus), .q(v1600obus), .dec(dec[1600]));
wire [data_w*2-1:0] v1601ibus;
wire [temp_w*2-1:0] v1601obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1601 (.l(l[1601*data_w +:data_w]), .r(v1601ibus), .q(v1601obus), .dec(dec[1601]));
wire [data_w*2-1:0] v1602ibus;
wire [temp_w*2-1:0] v1602obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1602 (.l(l[1602*data_w +:data_w]), .r(v1602ibus), .q(v1602obus), .dec(dec[1602]));
wire [data_w*2-1:0] v1603ibus;
wire [temp_w*2-1:0] v1603obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1603 (.l(l[1603*data_w +:data_w]), .r(v1603ibus), .q(v1603obus), .dec(dec[1603]));
wire [data_w*2-1:0] v1604ibus;
wire [temp_w*2-1:0] v1604obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1604 (.l(l[1604*data_w +:data_w]), .r(v1604ibus), .q(v1604obus), .dec(dec[1604]));
wire [data_w*2-1:0] v1605ibus;
wire [temp_w*2-1:0] v1605obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1605 (.l(l[1605*data_w +:data_w]), .r(v1605ibus), .q(v1605obus), .dec(dec[1605]));
wire [data_w*2-1:0] v1606ibus;
wire [temp_w*2-1:0] v1606obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1606 (.l(l[1606*data_w +:data_w]), .r(v1606ibus), .q(v1606obus), .dec(dec[1606]));
wire [data_w*2-1:0] v1607ibus;
wire [temp_w*2-1:0] v1607obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1607 (.l(l[1607*data_w +:data_w]), .r(v1607ibus), .q(v1607obus), .dec(dec[1607]));
wire [data_w*2-1:0] v1608ibus;
wire [temp_w*2-1:0] v1608obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1608 (.l(l[1608*data_w +:data_w]), .r(v1608ibus), .q(v1608obus), .dec(dec[1608]));
wire [data_w*2-1:0] v1609ibus;
wire [temp_w*2-1:0] v1609obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1609 (.l(l[1609*data_w +:data_w]), .r(v1609ibus), .q(v1609obus), .dec(dec[1609]));
wire [data_w*2-1:0] v1610ibus;
wire [temp_w*2-1:0] v1610obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1610 (.l(l[1610*data_w +:data_w]), .r(v1610ibus), .q(v1610obus), .dec(dec[1610]));
wire [data_w*2-1:0] v1611ibus;
wire [temp_w*2-1:0] v1611obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1611 (.l(l[1611*data_w +:data_w]), .r(v1611ibus), .q(v1611obus), .dec(dec[1611]));
wire [data_w*2-1:0] v1612ibus;
wire [temp_w*2-1:0] v1612obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1612 (.l(l[1612*data_w +:data_w]), .r(v1612ibus), .q(v1612obus), .dec(dec[1612]));
wire [data_w*2-1:0] v1613ibus;
wire [temp_w*2-1:0] v1613obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1613 (.l(l[1613*data_w +:data_w]), .r(v1613ibus), .q(v1613obus), .dec(dec[1613]));
wire [data_w*2-1:0] v1614ibus;
wire [temp_w*2-1:0] v1614obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1614 (.l(l[1614*data_w +:data_w]), .r(v1614ibus), .q(v1614obus), .dec(dec[1614]));
wire [data_w*2-1:0] v1615ibus;
wire [temp_w*2-1:0] v1615obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1615 (.l(l[1615*data_w +:data_w]), .r(v1615ibus), .q(v1615obus), .dec(dec[1615]));
wire [data_w*2-1:0] v1616ibus;
wire [temp_w*2-1:0] v1616obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1616 (.l(l[1616*data_w +:data_w]), .r(v1616ibus), .q(v1616obus), .dec(dec[1616]));
wire [data_w*2-1:0] v1617ibus;
wire [temp_w*2-1:0] v1617obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1617 (.l(l[1617*data_w +:data_w]), .r(v1617ibus), .q(v1617obus), .dec(dec[1617]));
wire [data_w*2-1:0] v1618ibus;
wire [temp_w*2-1:0] v1618obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1618 (.l(l[1618*data_w +:data_w]), .r(v1618ibus), .q(v1618obus), .dec(dec[1618]));
wire [data_w*2-1:0] v1619ibus;
wire [temp_w*2-1:0] v1619obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1619 (.l(l[1619*data_w +:data_w]), .r(v1619ibus), .q(v1619obus), .dec(dec[1619]));
wire [data_w*2-1:0] v1620ibus;
wire [temp_w*2-1:0] v1620obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1620 (.l(l[1620*data_w +:data_w]), .r(v1620ibus), .q(v1620obus), .dec(dec[1620]));
wire [data_w*2-1:0] v1621ibus;
wire [temp_w*2-1:0] v1621obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1621 (.l(l[1621*data_w +:data_w]), .r(v1621ibus), .q(v1621obus), .dec(dec[1621]));
wire [data_w*2-1:0] v1622ibus;
wire [temp_w*2-1:0] v1622obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1622 (.l(l[1622*data_w +:data_w]), .r(v1622ibus), .q(v1622obus), .dec(dec[1622]));
wire [data_w*2-1:0] v1623ibus;
wire [temp_w*2-1:0] v1623obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1623 (.l(l[1623*data_w +:data_w]), .r(v1623ibus), .q(v1623obus), .dec(dec[1623]));
wire [data_w*2-1:0] v1624ibus;
wire [temp_w*2-1:0] v1624obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1624 (.l(l[1624*data_w +:data_w]), .r(v1624ibus), .q(v1624obus), .dec(dec[1624]));
wire [data_w*2-1:0] v1625ibus;
wire [temp_w*2-1:0] v1625obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1625 (.l(l[1625*data_w +:data_w]), .r(v1625ibus), .q(v1625obus), .dec(dec[1625]));
wire [data_w*2-1:0] v1626ibus;
wire [temp_w*2-1:0] v1626obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1626 (.l(l[1626*data_w +:data_w]), .r(v1626ibus), .q(v1626obus), .dec(dec[1626]));
wire [data_w*2-1:0] v1627ibus;
wire [temp_w*2-1:0] v1627obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1627 (.l(l[1627*data_w +:data_w]), .r(v1627ibus), .q(v1627obus), .dec(dec[1627]));
wire [data_w*2-1:0] v1628ibus;
wire [temp_w*2-1:0] v1628obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1628 (.l(l[1628*data_w +:data_w]), .r(v1628ibus), .q(v1628obus), .dec(dec[1628]));
wire [data_w*2-1:0] v1629ibus;
wire [temp_w*2-1:0] v1629obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1629 (.l(l[1629*data_w +:data_w]), .r(v1629ibus), .q(v1629obus), .dec(dec[1629]));
wire [data_w*2-1:0] v1630ibus;
wire [temp_w*2-1:0] v1630obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1630 (.l(l[1630*data_w +:data_w]), .r(v1630ibus), .q(v1630obus), .dec(dec[1630]));
wire [data_w*2-1:0] v1631ibus;
wire [temp_w*2-1:0] v1631obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1631 (.l(l[1631*data_w +:data_w]), .r(v1631ibus), .q(v1631obus), .dec(dec[1631]));
wire [data_w*2-1:0] v1632ibus;
wire [temp_w*2-1:0] v1632obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1632 (.l(l[1632*data_w +:data_w]), .r(v1632ibus), .q(v1632obus), .dec(dec[1632]));
wire [data_w*2-1:0] v1633ibus;
wire [temp_w*2-1:0] v1633obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1633 (.l(l[1633*data_w +:data_w]), .r(v1633ibus), .q(v1633obus), .dec(dec[1633]));
wire [data_w*2-1:0] v1634ibus;
wire [temp_w*2-1:0] v1634obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1634 (.l(l[1634*data_w +:data_w]), .r(v1634ibus), .q(v1634obus), .dec(dec[1634]));
wire [data_w*2-1:0] v1635ibus;
wire [temp_w*2-1:0] v1635obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1635 (.l(l[1635*data_w +:data_w]), .r(v1635ibus), .q(v1635obus), .dec(dec[1635]));
wire [data_w*2-1:0] v1636ibus;
wire [temp_w*2-1:0] v1636obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1636 (.l(l[1636*data_w +:data_w]), .r(v1636ibus), .q(v1636obus), .dec(dec[1636]));
wire [data_w*2-1:0] v1637ibus;
wire [temp_w*2-1:0] v1637obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1637 (.l(l[1637*data_w +:data_w]), .r(v1637ibus), .q(v1637obus), .dec(dec[1637]));
wire [data_w*2-1:0] v1638ibus;
wire [temp_w*2-1:0] v1638obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1638 (.l(l[1638*data_w +:data_w]), .r(v1638ibus), .q(v1638obus), .dec(dec[1638]));
wire [data_w*2-1:0] v1639ibus;
wire [temp_w*2-1:0] v1639obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1639 (.l(l[1639*data_w +:data_w]), .r(v1639ibus), .q(v1639obus), .dec(dec[1639]));
wire [data_w*2-1:0] v1640ibus;
wire [temp_w*2-1:0] v1640obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1640 (.l(l[1640*data_w +:data_w]), .r(v1640ibus), .q(v1640obus), .dec(dec[1640]));
wire [data_w*2-1:0] v1641ibus;
wire [temp_w*2-1:0] v1641obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1641 (.l(l[1641*data_w +:data_w]), .r(v1641ibus), .q(v1641obus), .dec(dec[1641]));
wire [data_w*2-1:0] v1642ibus;
wire [temp_w*2-1:0] v1642obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1642 (.l(l[1642*data_w +:data_w]), .r(v1642ibus), .q(v1642obus), .dec(dec[1642]));
wire [data_w*2-1:0] v1643ibus;
wire [temp_w*2-1:0] v1643obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1643 (.l(l[1643*data_w +:data_w]), .r(v1643ibus), .q(v1643obus), .dec(dec[1643]));
wire [data_w*2-1:0] v1644ibus;
wire [temp_w*2-1:0] v1644obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1644 (.l(l[1644*data_w +:data_w]), .r(v1644ibus), .q(v1644obus), .dec(dec[1644]));
wire [data_w*2-1:0] v1645ibus;
wire [temp_w*2-1:0] v1645obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1645 (.l(l[1645*data_w +:data_w]), .r(v1645ibus), .q(v1645obus), .dec(dec[1645]));
wire [data_w*2-1:0] v1646ibus;
wire [temp_w*2-1:0] v1646obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1646 (.l(l[1646*data_w +:data_w]), .r(v1646ibus), .q(v1646obus), .dec(dec[1646]));
wire [data_w*2-1:0] v1647ibus;
wire [temp_w*2-1:0] v1647obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1647 (.l(l[1647*data_w +:data_w]), .r(v1647ibus), .q(v1647obus), .dec(dec[1647]));
wire [data_w*2-1:0] v1648ibus;
wire [temp_w*2-1:0] v1648obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1648 (.l(l[1648*data_w +:data_w]), .r(v1648ibus), .q(v1648obus), .dec(dec[1648]));
wire [data_w*2-1:0] v1649ibus;
wire [temp_w*2-1:0] v1649obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1649 (.l(l[1649*data_w +:data_w]), .r(v1649ibus), .q(v1649obus), .dec(dec[1649]));
wire [data_w*2-1:0] v1650ibus;
wire [temp_w*2-1:0] v1650obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1650 (.l(l[1650*data_w +:data_w]), .r(v1650ibus), .q(v1650obus), .dec(dec[1650]));
wire [data_w*2-1:0] v1651ibus;
wire [temp_w*2-1:0] v1651obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1651 (.l(l[1651*data_w +:data_w]), .r(v1651ibus), .q(v1651obus), .dec(dec[1651]));
wire [data_w*2-1:0] v1652ibus;
wire [temp_w*2-1:0] v1652obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1652 (.l(l[1652*data_w +:data_w]), .r(v1652ibus), .q(v1652obus), .dec(dec[1652]));
wire [data_w*2-1:0] v1653ibus;
wire [temp_w*2-1:0] v1653obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1653 (.l(l[1653*data_w +:data_w]), .r(v1653ibus), .q(v1653obus), .dec(dec[1653]));
wire [data_w*2-1:0] v1654ibus;
wire [temp_w*2-1:0] v1654obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1654 (.l(l[1654*data_w +:data_w]), .r(v1654ibus), .q(v1654obus), .dec(dec[1654]));
wire [data_w*2-1:0] v1655ibus;
wire [temp_w*2-1:0] v1655obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1655 (.l(l[1655*data_w +:data_w]), .r(v1655ibus), .q(v1655obus), .dec(dec[1655]));
wire [data_w*2-1:0] v1656ibus;
wire [temp_w*2-1:0] v1656obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1656 (.l(l[1656*data_w +:data_w]), .r(v1656ibus), .q(v1656obus), .dec(dec[1656]));
wire [data_w*2-1:0] v1657ibus;
wire [temp_w*2-1:0] v1657obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1657 (.l(l[1657*data_w +:data_w]), .r(v1657ibus), .q(v1657obus), .dec(dec[1657]));
wire [data_w*2-1:0] v1658ibus;
wire [temp_w*2-1:0] v1658obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1658 (.l(l[1658*data_w +:data_w]), .r(v1658ibus), .q(v1658obus), .dec(dec[1658]));
wire [data_w*2-1:0] v1659ibus;
wire [temp_w*2-1:0] v1659obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1659 (.l(l[1659*data_w +:data_w]), .r(v1659ibus), .q(v1659obus), .dec(dec[1659]));
wire [data_w*2-1:0] v1660ibus;
wire [temp_w*2-1:0] v1660obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1660 (.l(l[1660*data_w +:data_w]), .r(v1660ibus), .q(v1660obus), .dec(dec[1660]));
wire [data_w*2-1:0] v1661ibus;
wire [temp_w*2-1:0] v1661obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1661 (.l(l[1661*data_w +:data_w]), .r(v1661ibus), .q(v1661obus), .dec(dec[1661]));
wire [data_w*2-1:0] v1662ibus;
wire [temp_w*2-1:0] v1662obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1662 (.l(l[1662*data_w +:data_w]), .r(v1662ibus), .q(v1662obus), .dec(dec[1662]));
wire [data_w*2-1:0] v1663ibus;
wire [temp_w*2-1:0] v1663obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1663 (.l(l[1663*data_w +:data_w]), .r(v1663ibus), .q(v1663obus), .dec(dec[1663]));
wire [data_w*2-1:0] v1664ibus;
wire [temp_w*2-1:0] v1664obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1664 (.l(l[1664*data_w +:data_w]), .r(v1664ibus), .q(v1664obus), .dec(dec[1664]));
wire [data_w*2-1:0] v1665ibus;
wire [temp_w*2-1:0] v1665obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1665 (.l(l[1665*data_w +:data_w]), .r(v1665ibus), .q(v1665obus), .dec(dec[1665]));
wire [data_w*2-1:0] v1666ibus;
wire [temp_w*2-1:0] v1666obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1666 (.l(l[1666*data_w +:data_w]), .r(v1666ibus), .q(v1666obus), .dec(dec[1666]));
wire [data_w*2-1:0] v1667ibus;
wire [temp_w*2-1:0] v1667obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1667 (.l(l[1667*data_w +:data_w]), .r(v1667ibus), .q(v1667obus), .dec(dec[1667]));
wire [data_w*2-1:0] v1668ibus;
wire [temp_w*2-1:0] v1668obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1668 (.l(l[1668*data_w +:data_w]), .r(v1668ibus), .q(v1668obus), .dec(dec[1668]));
wire [data_w*2-1:0] v1669ibus;
wire [temp_w*2-1:0] v1669obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1669 (.l(l[1669*data_w +:data_w]), .r(v1669ibus), .q(v1669obus), .dec(dec[1669]));
wire [data_w*2-1:0] v1670ibus;
wire [temp_w*2-1:0] v1670obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1670 (.l(l[1670*data_w +:data_w]), .r(v1670ibus), .q(v1670obus), .dec(dec[1670]));
wire [data_w*2-1:0] v1671ibus;
wire [temp_w*2-1:0] v1671obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1671 (.l(l[1671*data_w +:data_w]), .r(v1671ibus), .q(v1671obus), .dec(dec[1671]));
wire [data_w*2-1:0] v1672ibus;
wire [temp_w*2-1:0] v1672obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1672 (.l(l[1672*data_w +:data_w]), .r(v1672ibus), .q(v1672obus), .dec(dec[1672]));
wire [data_w*2-1:0] v1673ibus;
wire [temp_w*2-1:0] v1673obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1673 (.l(l[1673*data_w +:data_w]), .r(v1673ibus), .q(v1673obus), .dec(dec[1673]));
wire [data_w*2-1:0] v1674ibus;
wire [temp_w*2-1:0] v1674obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1674 (.l(l[1674*data_w +:data_w]), .r(v1674ibus), .q(v1674obus), .dec(dec[1674]));
wire [data_w*2-1:0] v1675ibus;
wire [temp_w*2-1:0] v1675obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1675 (.l(l[1675*data_w +:data_w]), .r(v1675ibus), .q(v1675obus), .dec(dec[1675]));
wire [data_w*2-1:0] v1676ibus;
wire [temp_w*2-1:0] v1676obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1676 (.l(l[1676*data_w +:data_w]), .r(v1676ibus), .q(v1676obus), .dec(dec[1676]));
wire [data_w*2-1:0] v1677ibus;
wire [temp_w*2-1:0] v1677obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1677 (.l(l[1677*data_w +:data_w]), .r(v1677ibus), .q(v1677obus), .dec(dec[1677]));
wire [data_w*2-1:0] v1678ibus;
wire [temp_w*2-1:0] v1678obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1678 (.l(l[1678*data_w +:data_w]), .r(v1678ibus), .q(v1678obus), .dec(dec[1678]));
wire [data_w*2-1:0] v1679ibus;
wire [temp_w*2-1:0] v1679obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1679 (.l(l[1679*data_w +:data_w]), .r(v1679ibus), .q(v1679obus), .dec(dec[1679]));
wire [data_w*2-1:0] v1680ibus;
wire [temp_w*2-1:0] v1680obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1680 (.l(l[1680*data_w +:data_w]), .r(v1680ibus), .q(v1680obus), .dec(dec[1680]));
wire [data_w*2-1:0] v1681ibus;
wire [temp_w*2-1:0] v1681obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1681 (.l(l[1681*data_w +:data_w]), .r(v1681ibus), .q(v1681obus), .dec(dec[1681]));
wire [data_w*2-1:0] v1682ibus;
wire [temp_w*2-1:0] v1682obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1682 (.l(l[1682*data_w +:data_w]), .r(v1682ibus), .q(v1682obus), .dec(dec[1682]));
wire [data_w*2-1:0] v1683ibus;
wire [temp_w*2-1:0] v1683obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1683 (.l(l[1683*data_w +:data_w]), .r(v1683ibus), .q(v1683obus), .dec(dec[1683]));
wire [data_w*2-1:0] v1684ibus;
wire [temp_w*2-1:0] v1684obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1684 (.l(l[1684*data_w +:data_w]), .r(v1684ibus), .q(v1684obus), .dec(dec[1684]));
wire [data_w*2-1:0] v1685ibus;
wire [temp_w*2-1:0] v1685obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1685 (.l(l[1685*data_w +:data_w]), .r(v1685ibus), .q(v1685obus), .dec(dec[1685]));
wire [data_w*2-1:0] v1686ibus;
wire [temp_w*2-1:0] v1686obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1686 (.l(l[1686*data_w +:data_w]), .r(v1686ibus), .q(v1686obus), .dec(dec[1686]));
wire [data_w*2-1:0] v1687ibus;
wire [temp_w*2-1:0] v1687obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1687 (.l(l[1687*data_w +:data_w]), .r(v1687ibus), .q(v1687obus), .dec(dec[1687]));
wire [data_w*2-1:0] v1688ibus;
wire [temp_w*2-1:0] v1688obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1688 (.l(l[1688*data_w +:data_w]), .r(v1688ibus), .q(v1688obus), .dec(dec[1688]));
wire [data_w*2-1:0] v1689ibus;
wire [temp_w*2-1:0] v1689obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1689 (.l(l[1689*data_w +:data_w]), .r(v1689ibus), .q(v1689obus), .dec(dec[1689]));
wire [data_w*2-1:0] v1690ibus;
wire [temp_w*2-1:0] v1690obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1690 (.l(l[1690*data_w +:data_w]), .r(v1690ibus), .q(v1690obus), .dec(dec[1690]));
wire [data_w*2-1:0] v1691ibus;
wire [temp_w*2-1:0] v1691obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1691 (.l(l[1691*data_w +:data_w]), .r(v1691ibus), .q(v1691obus), .dec(dec[1691]));
wire [data_w*2-1:0] v1692ibus;
wire [temp_w*2-1:0] v1692obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1692 (.l(l[1692*data_w +:data_w]), .r(v1692ibus), .q(v1692obus), .dec(dec[1692]));
wire [data_w*2-1:0] v1693ibus;
wire [temp_w*2-1:0] v1693obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1693 (.l(l[1693*data_w +:data_w]), .r(v1693ibus), .q(v1693obus), .dec(dec[1693]));
wire [data_w*2-1:0] v1694ibus;
wire [temp_w*2-1:0] v1694obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1694 (.l(l[1694*data_w +:data_w]), .r(v1694ibus), .q(v1694obus), .dec(dec[1694]));
wire [data_w*2-1:0] v1695ibus;
wire [temp_w*2-1:0] v1695obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1695 (.l(l[1695*data_w +:data_w]), .r(v1695ibus), .q(v1695obus), .dec(dec[1695]));
wire [data_w*2-1:0] v1696ibus;
wire [temp_w*2-1:0] v1696obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1696 (.l(l[1696*data_w +:data_w]), .r(v1696ibus), .q(v1696obus), .dec(dec[1696]));
wire [data_w*2-1:0] v1697ibus;
wire [temp_w*2-1:0] v1697obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1697 (.l(l[1697*data_w +:data_w]), .r(v1697ibus), .q(v1697obus), .dec(dec[1697]));
wire [data_w*2-1:0] v1698ibus;
wire [temp_w*2-1:0] v1698obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1698 (.l(l[1698*data_w +:data_w]), .r(v1698ibus), .q(v1698obus), .dec(dec[1698]));
wire [data_w*2-1:0] v1699ibus;
wire [temp_w*2-1:0] v1699obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1699 (.l(l[1699*data_w +:data_w]), .r(v1699ibus), .q(v1699obus), .dec(dec[1699]));
wire [data_w*2-1:0] v1700ibus;
wire [temp_w*2-1:0] v1700obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1700 (.l(l[1700*data_w +:data_w]), .r(v1700ibus), .q(v1700obus), .dec(dec[1700]));
wire [data_w*2-1:0] v1701ibus;
wire [temp_w*2-1:0] v1701obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1701 (.l(l[1701*data_w +:data_w]), .r(v1701ibus), .q(v1701obus), .dec(dec[1701]));
wire [data_w*2-1:0] v1702ibus;
wire [temp_w*2-1:0] v1702obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1702 (.l(l[1702*data_w +:data_w]), .r(v1702ibus), .q(v1702obus), .dec(dec[1702]));
wire [data_w*2-1:0] v1703ibus;
wire [temp_w*2-1:0] v1703obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1703 (.l(l[1703*data_w +:data_w]), .r(v1703ibus), .q(v1703obus), .dec(dec[1703]));
wire [data_w*2-1:0] v1704ibus;
wire [temp_w*2-1:0] v1704obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1704 (.l(l[1704*data_w +:data_w]), .r(v1704ibus), .q(v1704obus), .dec(dec[1704]));
wire [data_w*2-1:0] v1705ibus;
wire [temp_w*2-1:0] v1705obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1705 (.l(l[1705*data_w +:data_w]), .r(v1705ibus), .q(v1705obus), .dec(dec[1705]));
wire [data_w*2-1:0] v1706ibus;
wire [temp_w*2-1:0] v1706obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1706 (.l(l[1706*data_w +:data_w]), .r(v1706ibus), .q(v1706obus), .dec(dec[1706]));
wire [data_w*2-1:0] v1707ibus;
wire [temp_w*2-1:0] v1707obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1707 (.l(l[1707*data_w +:data_w]), .r(v1707ibus), .q(v1707obus), .dec(dec[1707]));
wire [data_w*2-1:0] v1708ibus;
wire [temp_w*2-1:0] v1708obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1708 (.l(l[1708*data_w +:data_w]), .r(v1708ibus), .q(v1708obus), .dec(dec[1708]));
wire [data_w*2-1:0] v1709ibus;
wire [temp_w*2-1:0] v1709obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1709 (.l(l[1709*data_w +:data_w]), .r(v1709ibus), .q(v1709obus), .dec(dec[1709]));
wire [data_w*2-1:0] v1710ibus;
wire [temp_w*2-1:0] v1710obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1710 (.l(l[1710*data_w +:data_w]), .r(v1710ibus), .q(v1710obus), .dec(dec[1710]));
wire [data_w*2-1:0] v1711ibus;
wire [temp_w*2-1:0] v1711obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1711 (.l(l[1711*data_w +:data_w]), .r(v1711ibus), .q(v1711obus), .dec(dec[1711]));
wire [data_w*2-1:0] v1712ibus;
wire [temp_w*2-1:0] v1712obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1712 (.l(l[1712*data_w +:data_w]), .r(v1712ibus), .q(v1712obus), .dec(dec[1712]));
wire [data_w*2-1:0] v1713ibus;
wire [temp_w*2-1:0] v1713obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1713 (.l(l[1713*data_w +:data_w]), .r(v1713ibus), .q(v1713obus), .dec(dec[1713]));
wire [data_w*2-1:0] v1714ibus;
wire [temp_w*2-1:0] v1714obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1714 (.l(l[1714*data_w +:data_w]), .r(v1714ibus), .q(v1714obus), .dec(dec[1714]));
wire [data_w*2-1:0] v1715ibus;
wire [temp_w*2-1:0] v1715obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1715 (.l(l[1715*data_w +:data_w]), .r(v1715ibus), .q(v1715obus), .dec(dec[1715]));
wire [data_w*2-1:0] v1716ibus;
wire [temp_w*2-1:0] v1716obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1716 (.l(l[1716*data_w +:data_w]), .r(v1716ibus), .q(v1716obus), .dec(dec[1716]));
wire [data_w*2-1:0] v1717ibus;
wire [temp_w*2-1:0] v1717obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1717 (.l(l[1717*data_w +:data_w]), .r(v1717ibus), .q(v1717obus), .dec(dec[1717]));
wire [data_w*2-1:0] v1718ibus;
wire [temp_w*2-1:0] v1718obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1718 (.l(l[1718*data_w +:data_w]), .r(v1718ibus), .q(v1718obus), .dec(dec[1718]));
wire [data_w*2-1:0] v1719ibus;
wire [temp_w*2-1:0] v1719obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1719 (.l(l[1719*data_w +:data_w]), .r(v1719ibus), .q(v1719obus), .dec(dec[1719]));
wire [data_w*2-1:0] v1720ibus;
wire [temp_w*2-1:0] v1720obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1720 (.l(l[1720*data_w +:data_w]), .r(v1720ibus), .q(v1720obus), .dec(dec[1720]));
wire [data_w*2-1:0] v1721ibus;
wire [temp_w*2-1:0] v1721obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1721 (.l(l[1721*data_w +:data_w]), .r(v1721ibus), .q(v1721obus), .dec(dec[1721]));
wire [data_w*2-1:0] v1722ibus;
wire [temp_w*2-1:0] v1722obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1722 (.l(l[1722*data_w +:data_w]), .r(v1722ibus), .q(v1722obus), .dec(dec[1722]));
wire [data_w*2-1:0] v1723ibus;
wire [temp_w*2-1:0] v1723obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1723 (.l(l[1723*data_w +:data_w]), .r(v1723ibus), .q(v1723obus), .dec(dec[1723]));
wire [data_w*2-1:0] v1724ibus;
wire [temp_w*2-1:0] v1724obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1724 (.l(l[1724*data_w +:data_w]), .r(v1724ibus), .q(v1724obus), .dec(dec[1724]));
wire [data_w*2-1:0] v1725ibus;
wire [temp_w*2-1:0] v1725obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1725 (.l(l[1725*data_w +:data_w]), .r(v1725ibus), .q(v1725obus), .dec(dec[1725]));
wire [data_w*2-1:0] v1726ibus;
wire [temp_w*2-1:0] v1726obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1726 (.l(l[1726*data_w +:data_w]), .r(v1726ibus), .q(v1726obus), .dec(dec[1726]));
wire [data_w*2-1:0] v1727ibus;
wire [temp_w*2-1:0] v1727obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1727 (.l(l[1727*data_w +:data_w]), .r(v1727ibus), .q(v1727obus), .dec(dec[1727]));
wire [data_w*2-1:0] v1728ibus;
wire [temp_w*2-1:0] v1728obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1728 (.l(l[1728*data_w +:data_w]), .r(v1728ibus), .q(v1728obus), .dec(dec[1728]));
wire [data_w*2-1:0] v1729ibus;
wire [temp_w*2-1:0] v1729obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1729 (.l(l[1729*data_w +:data_w]), .r(v1729ibus), .q(v1729obus), .dec(dec[1729]));
wire [data_w*2-1:0] v1730ibus;
wire [temp_w*2-1:0] v1730obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1730 (.l(l[1730*data_w +:data_w]), .r(v1730ibus), .q(v1730obus), .dec(dec[1730]));
wire [data_w*2-1:0] v1731ibus;
wire [temp_w*2-1:0] v1731obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1731 (.l(l[1731*data_w +:data_w]), .r(v1731ibus), .q(v1731obus), .dec(dec[1731]));
wire [data_w*2-1:0] v1732ibus;
wire [temp_w*2-1:0] v1732obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1732 (.l(l[1732*data_w +:data_w]), .r(v1732ibus), .q(v1732obus), .dec(dec[1732]));
wire [data_w*2-1:0] v1733ibus;
wire [temp_w*2-1:0] v1733obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1733 (.l(l[1733*data_w +:data_w]), .r(v1733ibus), .q(v1733obus), .dec(dec[1733]));
wire [data_w*2-1:0] v1734ibus;
wire [temp_w*2-1:0] v1734obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1734 (.l(l[1734*data_w +:data_w]), .r(v1734ibus), .q(v1734obus), .dec(dec[1734]));
wire [data_w*2-1:0] v1735ibus;
wire [temp_w*2-1:0] v1735obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1735 (.l(l[1735*data_w +:data_w]), .r(v1735ibus), .q(v1735obus), .dec(dec[1735]));
wire [data_w*2-1:0] v1736ibus;
wire [temp_w*2-1:0] v1736obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1736 (.l(l[1736*data_w +:data_w]), .r(v1736ibus), .q(v1736obus), .dec(dec[1736]));
wire [data_w*2-1:0] v1737ibus;
wire [temp_w*2-1:0] v1737obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1737 (.l(l[1737*data_w +:data_w]), .r(v1737ibus), .q(v1737obus), .dec(dec[1737]));
wire [data_w*2-1:0] v1738ibus;
wire [temp_w*2-1:0] v1738obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1738 (.l(l[1738*data_w +:data_w]), .r(v1738ibus), .q(v1738obus), .dec(dec[1738]));
wire [data_w*2-1:0] v1739ibus;
wire [temp_w*2-1:0] v1739obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1739 (.l(l[1739*data_w +:data_w]), .r(v1739ibus), .q(v1739obus), .dec(dec[1739]));
wire [data_w*2-1:0] v1740ibus;
wire [temp_w*2-1:0] v1740obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1740 (.l(l[1740*data_w +:data_w]), .r(v1740ibus), .q(v1740obus), .dec(dec[1740]));
wire [data_w*2-1:0] v1741ibus;
wire [temp_w*2-1:0] v1741obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1741 (.l(l[1741*data_w +:data_w]), .r(v1741ibus), .q(v1741obus), .dec(dec[1741]));
wire [data_w*2-1:0] v1742ibus;
wire [temp_w*2-1:0] v1742obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1742 (.l(l[1742*data_w +:data_w]), .r(v1742ibus), .q(v1742obus), .dec(dec[1742]));
wire [data_w*2-1:0] v1743ibus;
wire [temp_w*2-1:0] v1743obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1743 (.l(l[1743*data_w +:data_w]), .r(v1743ibus), .q(v1743obus), .dec(dec[1743]));
wire [data_w*2-1:0] v1744ibus;
wire [temp_w*2-1:0] v1744obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1744 (.l(l[1744*data_w +:data_w]), .r(v1744ibus), .q(v1744obus), .dec(dec[1744]));
wire [data_w*2-1:0] v1745ibus;
wire [temp_w*2-1:0] v1745obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1745 (.l(l[1745*data_w +:data_w]), .r(v1745ibus), .q(v1745obus), .dec(dec[1745]));
wire [data_w*2-1:0] v1746ibus;
wire [temp_w*2-1:0] v1746obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1746 (.l(l[1746*data_w +:data_w]), .r(v1746ibus), .q(v1746obus), .dec(dec[1746]));
wire [data_w*2-1:0] v1747ibus;
wire [temp_w*2-1:0] v1747obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1747 (.l(l[1747*data_w +:data_w]), .r(v1747ibus), .q(v1747obus), .dec(dec[1747]));
wire [data_w*2-1:0] v1748ibus;
wire [temp_w*2-1:0] v1748obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1748 (.l(l[1748*data_w +:data_w]), .r(v1748ibus), .q(v1748obus), .dec(dec[1748]));
wire [data_w*2-1:0] v1749ibus;
wire [temp_w*2-1:0] v1749obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1749 (.l(l[1749*data_w +:data_w]), .r(v1749ibus), .q(v1749obus), .dec(dec[1749]));
wire [data_w*2-1:0] v1750ibus;
wire [temp_w*2-1:0] v1750obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1750 (.l(l[1750*data_w +:data_w]), .r(v1750ibus), .q(v1750obus), .dec(dec[1750]));
wire [data_w*2-1:0] v1751ibus;
wire [temp_w*2-1:0] v1751obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1751 (.l(l[1751*data_w +:data_w]), .r(v1751ibus), .q(v1751obus), .dec(dec[1751]));
wire [data_w*2-1:0] v1752ibus;
wire [temp_w*2-1:0] v1752obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1752 (.l(l[1752*data_w +:data_w]), .r(v1752ibus), .q(v1752obus), .dec(dec[1752]));
wire [data_w*2-1:0] v1753ibus;
wire [temp_w*2-1:0] v1753obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1753 (.l(l[1753*data_w +:data_w]), .r(v1753ibus), .q(v1753obus), .dec(dec[1753]));
wire [data_w*2-1:0] v1754ibus;
wire [temp_w*2-1:0] v1754obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1754 (.l(l[1754*data_w +:data_w]), .r(v1754ibus), .q(v1754obus), .dec(dec[1754]));
wire [data_w*2-1:0] v1755ibus;
wire [temp_w*2-1:0] v1755obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1755 (.l(l[1755*data_w +:data_w]), .r(v1755ibus), .q(v1755obus), .dec(dec[1755]));
wire [data_w*2-1:0] v1756ibus;
wire [temp_w*2-1:0] v1756obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1756 (.l(l[1756*data_w +:data_w]), .r(v1756ibus), .q(v1756obus), .dec(dec[1756]));
wire [data_w*2-1:0] v1757ibus;
wire [temp_w*2-1:0] v1757obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1757 (.l(l[1757*data_w +:data_w]), .r(v1757ibus), .q(v1757obus), .dec(dec[1757]));
wire [data_w*2-1:0] v1758ibus;
wire [temp_w*2-1:0] v1758obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1758 (.l(l[1758*data_w +:data_w]), .r(v1758ibus), .q(v1758obus), .dec(dec[1758]));
wire [data_w*2-1:0] v1759ibus;
wire [temp_w*2-1:0] v1759obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1759 (.l(l[1759*data_w +:data_w]), .r(v1759ibus), .q(v1759obus), .dec(dec[1759]));
wire [data_w*2-1:0] v1760ibus;
wire [temp_w*2-1:0] v1760obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1760 (.l(l[1760*data_w +:data_w]), .r(v1760ibus), .q(v1760obus), .dec(dec[1760]));
wire [data_w*2-1:0] v1761ibus;
wire [temp_w*2-1:0] v1761obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1761 (.l(l[1761*data_w +:data_w]), .r(v1761ibus), .q(v1761obus), .dec(dec[1761]));
wire [data_w*2-1:0] v1762ibus;
wire [temp_w*2-1:0] v1762obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1762 (.l(l[1762*data_w +:data_w]), .r(v1762ibus), .q(v1762obus), .dec(dec[1762]));
wire [data_w*2-1:0] v1763ibus;
wire [temp_w*2-1:0] v1763obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1763 (.l(l[1763*data_w +:data_w]), .r(v1763ibus), .q(v1763obus), .dec(dec[1763]));
wire [data_w*2-1:0] v1764ibus;
wire [temp_w*2-1:0] v1764obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1764 (.l(l[1764*data_w +:data_w]), .r(v1764ibus), .q(v1764obus), .dec(dec[1764]));
wire [data_w*2-1:0] v1765ibus;
wire [temp_w*2-1:0] v1765obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1765 (.l(l[1765*data_w +:data_w]), .r(v1765ibus), .q(v1765obus), .dec(dec[1765]));
wire [data_w*2-1:0] v1766ibus;
wire [temp_w*2-1:0] v1766obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1766 (.l(l[1766*data_w +:data_w]), .r(v1766ibus), .q(v1766obus), .dec(dec[1766]));
wire [data_w*2-1:0] v1767ibus;
wire [temp_w*2-1:0] v1767obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1767 (.l(l[1767*data_w +:data_w]), .r(v1767ibus), .q(v1767obus), .dec(dec[1767]));
wire [data_w*2-1:0] v1768ibus;
wire [temp_w*2-1:0] v1768obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1768 (.l(l[1768*data_w +:data_w]), .r(v1768ibus), .q(v1768obus), .dec(dec[1768]));
wire [data_w*2-1:0] v1769ibus;
wire [temp_w*2-1:0] v1769obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1769 (.l(l[1769*data_w +:data_w]), .r(v1769ibus), .q(v1769obus), .dec(dec[1769]));
wire [data_w*2-1:0] v1770ibus;
wire [temp_w*2-1:0] v1770obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1770 (.l(l[1770*data_w +:data_w]), .r(v1770ibus), .q(v1770obus), .dec(dec[1770]));
wire [data_w*2-1:0] v1771ibus;
wire [temp_w*2-1:0] v1771obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1771 (.l(l[1771*data_w +:data_w]), .r(v1771ibus), .q(v1771obus), .dec(dec[1771]));
wire [data_w*2-1:0] v1772ibus;
wire [temp_w*2-1:0] v1772obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1772 (.l(l[1772*data_w +:data_w]), .r(v1772ibus), .q(v1772obus), .dec(dec[1772]));
wire [data_w*2-1:0] v1773ibus;
wire [temp_w*2-1:0] v1773obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1773 (.l(l[1773*data_w +:data_w]), .r(v1773ibus), .q(v1773obus), .dec(dec[1773]));
wire [data_w*2-1:0] v1774ibus;
wire [temp_w*2-1:0] v1774obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1774 (.l(l[1774*data_w +:data_w]), .r(v1774ibus), .q(v1774obus), .dec(dec[1774]));
wire [data_w*2-1:0] v1775ibus;
wire [temp_w*2-1:0] v1775obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1775 (.l(l[1775*data_w +:data_w]), .r(v1775ibus), .q(v1775obus), .dec(dec[1775]));
wire [data_w*2-1:0] v1776ibus;
wire [temp_w*2-1:0] v1776obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1776 (.l(l[1776*data_w +:data_w]), .r(v1776ibus), .q(v1776obus), .dec(dec[1776]));
wire [data_w*2-1:0] v1777ibus;
wire [temp_w*2-1:0] v1777obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1777 (.l(l[1777*data_w +:data_w]), .r(v1777ibus), .q(v1777obus), .dec(dec[1777]));
wire [data_w*2-1:0] v1778ibus;
wire [temp_w*2-1:0] v1778obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1778 (.l(l[1778*data_w +:data_w]), .r(v1778ibus), .q(v1778obus), .dec(dec[1778]));
wire [data_w*2-1:0] v1779ibus;
wire [temp_w*2-1:0] v1779obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1779 (.l(l[1779*data_w +:data_w]), .r(v1779ibus), .q(v1779obus), .dec(dec[1779]));
wire [data_w*2-1:0] v1780ibus;
wire [temp_w*2-1:0] v1780obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1780 (.l(l[1780*data_w +:data_w]), .r(v1780ibus), .q(v1780obus), .dec(dec[1780]));
wire [data_w*2-1:0] v1781ibus;
wire [temp_w*2-1:0] v1781obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1781 (.l(l[1781*data_w +:data_w]), .r(v1781ibus), .q(v1781obus), .dec(dec[1781]));
wire [data_w*2-1:0] v1782ibus;
wire [temp_w*2-1:0] v1782obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1782 (.l(l[1782*data_w +:data_w]), .r(v1782ibus), .q(v1782obus), .dec(dec[1782]));
wire [data_w*2-1:0] v1783ibus;
wire [temp_w*2-1:0] v1783obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1783 (.l(l[1783*data_w +:data_w]), .r(v1783ibus), .q(v1783obus), .dec(dec[1783]));
wire [data_w*2-1:0] v1784ibus;
wire [temp_w*2-1:0] v1784obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1784 (.l(l[1784*data_w +:data_w]), .r(v1784ibus), .q(v1784obus), .dec(dec[1784]));
wire [data_w*2-1:0] v1785ibus;
wire [temp_w*2-1:0] v1785obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1785 (.l(l[1785*data_w +:data_w]), .r(v1785ibus), .q(v1785obus), .dec(dec[1785]));
wire [data_w*2-1:0] v1786ibus;
wire [temp_w*2-1:0] v1786obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1786 (.l(l[1786*data_w +:data_w]), .r(v1786ibus), .q(v1786obus), .dec(dec[1786]));
wire [data_w*2-1:0] v1787ibus;
wire [temp_w*2-1:0] v1787obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1787 (.l(l[1787*data_w +:data_w]), .r(v1787ibus), .q(v1787obus), .dec(dec[1787]));
wire [data_w*2-1:0] v1788ibus;
wire [temp_w*2-1:0] v1788obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1788 (.l(l[1788*data_w +:data_w]), .r(v1788ibus), .q(v1788obus), .dec(dec[1788]));
wire [data_w*2-1:0] v1789ibus;
wire [temp_w*2-1:0] v1789obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1789 (.l(l[1789*data_w +:data_w]), .r(v1789ibus), .q(v1789obus), .dec(dec[1789]));
wire [data_w*2-1:0] v1790ibus;
wire [temp_w*2-1:0] v1790obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1790 (.l(l[1790*data_w +:data_w]), .r(v1790ibus), .q(v1790obus), .dec(dec[1790]));
wire [data_w*2-1:0] v1791ibus;
wire [temp_w*2-1:0] v1791obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1791 (.l(l[1791*data_w +:data_w]), .r(v1791ibus), .q(v1791obus), .dec(dec[1791]));
wire [data_w*2-1:0] v1792ibus;
wire [temp_w*2-1:0] v1792obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1792 (.l(l[1792*data_w +:data_w]), .r(v1792ibus), .q(v1792obus), .dec(dec[1792]));
wire [data_w*2-1:0] v1793ibus;
wire [temp_w*2-1:0] v1793obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1793 (.l(l[1793*data_w +:data_w]), .r(v1793ibus), .q(v1793obus), .dec(dec[1793]));
wire [data_w*2-1:0] v1794ibus;
wire [temp_w*2-1:0] v1794obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1794 (.l(l[1794*data_w +:data_w]), .r(v1794ibus), .q(v1794obus), .dec(dec[1794]));
wire [data_w*2-1:0] v1795ibus;
wire [temp_w*2-1:0] v1795obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1795 (.l(l[1795*data_w +:data_w]), .r(v1795ibus), .q(v1795obus), .dec(dec[1795]));
wire [data_w*2-1:0] v1796ibus;
wire [temp_w*2-1:0] v1796obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1796 (.l(l[1796*data_w +:data_w]), .r(v1796ibus), .q(v1796obus), .dec(dec[1796]));
wire [data_w*2-1:0] v1797ibus;
wire [temp_w*2-1:0] v1797obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1797 (.l(l[1797*data_w +:data_w]), .r(v1797ibus), .q(v1797obus), .dec(dec[1797]));
wire [data_w*2-1:0] v1798ibus;
wire [temp_w*2-1:0] v1798obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1798 (.l(l[1798*data_w +:data_w]), .r(v1798ibus), .q(v1798obus), .dec(dec[1798]));
wire [data_w*2-1:0] v1799ibus;
wire [temp_w*2-1:0] v1799obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1799 (.l(l[1799*data_w +:data_w]), .r(v1799ibus), .q(v1799obus), .dec(dec[1799]));
wire [data_w*2-1:0] v1800ibus;
wire [temp_w*2-1:0] v1800obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1800 (.l(l[1800*data_w +:data_w]), .r(v1800ibus), .q(v1800obus), .dec(dec[1800]));
wire [data_w*2-1:0] v1801ibus;
wire [temp_w*2-1:0] v1801obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1801 (.l(l[1801*data_w +:data_w]), .r(v1801ibus), .q(v1801obus), .dec(dec[1801]));
wire [data_w*2-1:0] v1802ibus;
wire [temp_w*2-1:0] v1802obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1802 (.l(l[1802*data_w +:data_w]), .r(v1802ibus), .q(v1802obus), .dec(dec[1802]));
wire [data_w*2-1:0] v1803ibus;
wire [temp_w*2-1:0] v1803obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1803 (.l(l[1803*data_w +:data_w]), .r(v1803ibus), .q(v1803obus), .dec(dec[1803]));
wire [data_w*2-1:0] v1804ibus;
wire [temp_w*2-1:0] v1804obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1804 (.l(l[1804*data_w +:data_w]), .r(v1804ibus), .q(v1804obus), .dec(dec[1804]));
wire [data_w*2-1:0] v1805ibus;
wire [temp_w*2-1:0] v1805obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1805 (.l(l[1805*data_w +:data_w]), .r(v1805ibus), .q(v1805obus), .dec(dec[1805]));
wire [data_w*2-1:0] v1806ibus;
wire [temp_w*2-1:0] v1806obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1806 (.l(l[1806*data_w +:data_w]), .r(v1806ibus), .q(v1806obus), .dec(dec[1806]));
wire [data_w*2-1:0] v1807ibus;
wire [temp_w*2-1:0] v1807obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1807 (.l(l[1807*data_w +:data_w]), .r(v1807ibus), .q(v1807obus), .dec(dec[1807]));
wire [data_w*2-1:0] v1808ibus;
wire [temp_w*2-1:0] v1808obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1808 (.l(l[1808*data_w +:data_w]), .r(v1808ibus), .q(v1808obus), .dec(dec[1808]));
wire [data_w*2-1:0] v1809ibus;
wire [temp_w*2-1:0] v1809obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1809 (.l(l[1809*data_w +:data_w]), .r(v1809ibus), .q(v1809obus), .dec(dec[1809]));
wire [data_w*2-1:0] v1810ibus;
wire [temp_w*2-1:0] v1810obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1810 (.l(l[1810*data_w +:data_w]), .r(v1810ibus), .q(v1810obus), .dec(dec[1810]));
wire [data_w*2-1:0] v1811ibus;
wire [temp_w*2-1:0] v1811obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1811 (.l(l[1811*data_w +:data_w]), .r(v1811ibus), .q(v1811obus), .dec(dec[1811]));
wire [data_w*2-1:0] v1812ibus;
wire [temp_w*2-1:0] v1812obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1812 (.l(l[1812*data_w +:data_w]), .r(v1812ibus), .q(v1812obus), .dec(dec[1812]));
wire [data_w*2-1:0] v1813ibus;
wire [temp_w*2-1:0] v1813obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1813 (.l(l[1813*data_w +:data_w]), .r(v1813ibus), .q(v1813obus), .dec(dec[1813]));
wire [data_w*2-1:0] v1814ibus;
wire [temp_w*2-1:0] v1814obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1814 (.l(l[1814*data_w +:data_w]), .r(v1814ibus), .q(v1814obus), .dec(dec[1814]));
wire [data_w*2-1:0] v1815ibus;
wire [temp_w*2-1:0] v1815obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1815 (.l(l[1815*data_w +:data_w]), .r(v1815ibus), .q(v1815obus), .dec(dec[1815]));
wire [data_w*2-1:0] v1816ibus;
wire [temp_w*2-1:0] v1816obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1816 (.l(l[1816*data_w +:data_w]), .r(v1816ibus), .q(v1816obus), .dec(dec[1816]));
wire [data_w*2-1:0] v1817ibus;
wire [temp_w*2-1:0] v1817obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1817 (.l(l[1817*data_w +:data_w]), .r(v1817ibus), .q(v1817obus), .dec(dec[1817]));
wire [data_w*2-1:0] v1818ibus;
wire [temp_w*2-1:0] v1818obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1818 (.l(l[1818*data_w +:data_w]), .r(v1818ibus), .q(v1818obus), .dec(dec[1818]));
wire [data_w*2-1:0] v1819ibus;
wire [temp_w*2-1:0] v1819obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1819 (.l(l[1819*data_w +:data_w]), .r(v1819ibus), .q(v1819obus), .dec(dec[1819]));
wire [data_w*2-1:0] v1820ibus;
wire [temp_w*2-1:0] v1820obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1820 (.l(l[1820*data_w +:data_w]), .r(v1820ibus), .q(v1820obus), .dec(dec[1820]));
wire [data_w*2-1:0] v1821ibus;
wire [temp_w*2-1:0] v1821obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1821 (.l(l[1821*data_w +:data_w]), .r(v1821ibus), .q(v1821obus), .dec(dec[1821]));
wire [data_w*2-1:0] v1822ibus;
wire [temp_w*2-1:0] v1822obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1822 (.l(l[1822*data_w +:data_w]), .r(v1822ibus), .q(v1822obus), .dec(dec[1822]));
wire [data_w*2-1:0] v1823ibus;
wire [temp_w*2-1:0] v1823obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1823 (.l(l[1823*data_w +:data_w]), .r(v1823ibus), .q(v1823obus), .dec(dec[1823]));
wire [data_w*2-1:0] v1824ibus;
wire [temp_w*2-1:0] v1824obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1824 (.l(l[1824*data_w +:data_w]), .r(v1824ibus), .q(v1824obus), .dec(dec[1824]));
wire [data_w*2-1:0] v1825ibus;
wire [temp_w*2-1:0] v1825obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1825 (.l(l[1825*data_w +:data_w]), .r(v1825ibus), .q(v1825obus), .dec(dec[1825]));
wire [data_w*2-1:0] v1826ibus;
wire [temp_w*2-1:0] v1826obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1826 (.l(l[1826*data_w +:data_w]), .r(v1826ibus), .q(v1826obus), .dec(dec[1826]));
wire [data_w*2-1:0] v1827ibus;
wire [temp_w*2-1:0] v1827obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1827 (.l(l[1827*data_w +:data_w]), .r(v1827ibus), .q(v1827obus), .dec(dec[1827]));
wire [data_w*2-1:0] v1828ibus;
wire [temp_w*2-1:0] v1828obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1828 (.l(l[1828*data_w +:data_w]), .r(v1828ibus), .q(v1828obus), .dec(dec[1828]));
wire [data_w*2-1:0] v1829ibus;
wire [temp_w*2-1:0] v1829obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1829 (.l(l[1829*data_w +:data_w]), .r(v1829ibus), .q(v1829obus), .dec(dec[1829]));
wire [data_w*2-1:0] v1830ibus;
wire [temp_w*2-1:0] v1830obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1830 (.l(l[1830*data_w +:data_w]), .r(v1830ibus), .q(v1830obus), .dec(dec[1830]));
wire [data_w*2-1:0] v1831ibus;
wire [temp_w*2-1:0] v1831obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1831 (.l(l[1831*data_w +:data_w]), .r(v1831ibus), .q(v1831obus), .dec(dec[1831]));
wire [data_w*2-1:0] v1832ibus;
wire [temp_w*2-1:0] v1832obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1832 (.l(l[1832*data_w +:data_w]), .r(v1832ibus), .q(v1832obus), .dec(dec[1832]));
wire [data_w*2-1:0] v1833ibus;
wire [temp_w*2-1:0] v1833obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1833 (.l(l[1833*data_w +:data_w]), .r(v1833ibus), .q(v1833obus), .dec(dec[1833]));
wire [data_w*2-1:0] v1834ibus;
wire [temp_w*2-1:0] v1834obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1834 (.l(l[1834*data_w +:data_w]), .r(v1834ibus), .q(v1834obus), .dec(dec[1834]));
wire [data_w*2-1:0] v1835ibus;
wire [temp_w*2-1:0] v1835obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1835 (.l(l[1835*data_w +:data_w]), .r(v1835ibus), .q(v1835obus), .dec(dec[1835]));
wire [data_w*2-1:0] v1836ibus;
wire [temp_w*2-1:0] v1836obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1836 (.l(l[1836*data_w +:data_w]), .r(v1836ibus), .q(v1836obus), .dec(dec[1836]));
wire [data_w*2-1:0] v1837ibus;
wire [temp_w*2-1:0] v1837obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1837 (.l(l[1837*data_w +:data_w]), .r(v1837ibus), .q(v1837obus), .dec(dec[1837]));
wire [data_w*2-1:0] v1838ibus;
wire [temp_w*2-1:0] v1838obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1838 (.l(l[1838*data_w +:data_w]), .r(v1838ibus), .q(v1838obus), .dec(dec[1838]));
wire [data_w*2-1:0] v1839ibus;
wire [temp_w*2-1:0] v1839obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1839 (.l(l[1839*data_w +:data_w]), .r(v1839ibus), .q(v1839obus), .dec(dec[1839]));
wire [data_w*2-1:0] v1840ibus;
wire [temp_w*2-1:0] v1840obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1840 (.l(l[1840*data_w +:data_w]), .r(v1840ibus), .q(v1840obus), .dec(dec[1840]));
wire [data_w*2-1:0] v1841ibus;
wire [temp_w*2-1:0] v1841obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1841 (.l(l[1841*data_w +:data_w]), .r(v1841ibus), .q(v1841obus), .dec(dec[1841]));
wire [data_w*2-1:0] v1842ibus;
wire [temp_w*2-1:0] v1842obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1842 (.l(l[1842*data_w +:data_w]), .r(v1842ibus), .q(v1842obus), .dec(dec[1842]));
wire [data_w*2-1:0] v1843ibus;
wire [temp_w*2-1:0] v1843obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1843 (.l(l[1843*data_w +:data_w]), .r(v1843ibus), .q(v1843obus), .dec(dec[1843]));
wire [data_w*2-1:0] v1844ibus;
wire [temp_w*2-1:0] v1844obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1844 (.l(l[1844*data_w +:data_w]), .r(v1844ibus), .q(v1844obus), .dec(dec[1844]));
wire [data_w*2-1:0] v1845ibus;
wire [temp_w*2-1:0] v1845obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1845 (.l(l[1845*data_w +:data_w]), .r(v1845ibus), .q(v1845obus), .dec(dec[1845]));
wire [data_w*2-1:0] v1846ibus;
wire [temp_w*2-1:0] v1846obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1846 (.l(l[1846*data_w +:data_w]), .r(v1846ibus), .q(v1846obus), .dec(dec[1846]));
wire [data_w*2-1:0] v1847ibus;
wire [temp_w*2-1:0] v1847obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1847 (.l(l[1847*data_w +:data_w]), .r(v1847ibus), .q(v1847obus), .dec(dec[1847]));
wire [data_w*2-1:0] v1848ibus;
wire [temp_w*2-1:0] v1848obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1848 (.l(l[1848*data_w +:data_w]), .r(v1848ibus), .q(v1848obus), .dec(dec[1848]));
wire [data_w*2-1:0] v1849ibus;
wire [temp_w*2-1:0] v1849obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1849 (.l(l[1849*data_w +:data_w]), .r(v1849ibus), .q(v1849obus), .dec(dec[1849]));
wire [data_w*2-1:0] v1850ibus;
wire [temp_w*2-1:0] v1850obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1850 (.l(l[1850*data_w +:data_w]), .r(v1850ibus), .q(v1850obus), .dec(dec[1850]));
wire [data_w*2-1:0] v1851ibus;
wire [temp_w*2-1:0] v1851obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1851 (.l(l[1851*data_w +:data_w]), .r(v1851ibus), .q(v1851obus), .dec(dec[1851]));
wire [data_w*2-1:0] v1852ibus;
wire [temp_w*2-1:0] v1852obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1852 (.l(l[1852*data_w +:data_w]), .r(v1852ibus), .q(v1852obus), .dec(dec[1852]));
wire [data_w*2-1:0] v1853ibus;
wire [temp_w*2-1:0] v1853obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1853 (.l(l[1853*data_w +:data_w]), .r(v1853ibus), .q(v1853obus), .dec(dec[1853]));
wire [data_w*2-1:0] v1854ibus;
wire [temp_w*2-1:0] v1854obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1854 (.l(l[1854*data_w +:data_w]), .r(v1854ibus), .q(v1854obus), .dec(dec[1854]));
wire [data_w*2-1:0] v1855ibus;
wire [temp_w*2-1:0] v1855obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1855 (.l(l[1855*data_w +:data_w]), .r(v1855ibus), .q(v1855obus), .dec(dec[1855]));
wire [data_w*2-1:0] v1856ibus;
wire [temp_w*2-1:0] v1856obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1856 (.l(l[1856*data_w +:data_w]), .r(v1856ibus), .q(v1856obus), .dec(dec[1856]));
wire [data_w*2-1:0] v1857ibus;
wire [temp_w*2-1:0] v1857obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1857 (.l(l[1857*data_w +:data_w]), .r(v1857ibus), .q(v1857obus), .dec(dec[1857]));
wire [data_w*2-1:0] v1858ibus;
wire [temp_w*2-1:0] v1858obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1858 (.l(l[1858*data_w +:data_w]), .r(v1858ibus), .q(v1858obus), .dec(dec[1858]));
wire [data_w*2-1:0] v1859ibus;
wire [temp_w*2-1:0] v1859obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1859 (.l(l[1859*data_w +:data_w]), .r(v1859ibus), .q(v1859obus), .dec(dec[1859]));
wire [data_w*2-1:0] v1860ibus;
wire [temp_w*2-1:0] v1860obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1860 (.l(l[1860*data_w +:data_w]), .r(v1860ibus), .q(v1860obus), .dec(dec[1860]));
wire [data_w*2-1:0] v1861ibus;
wire [temp_w*2-1:0] v1861obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1861 (.l(l[1861*data_w +:data_w]), .r(v1861ibus), .q(v1861obus), .dec(dec[1861]));
wire [data_w*2-1:0] v1862ibus;
wire [temp_w*2-1:0] v1862obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1862 (.l(l[1862*data_w +:data_w]), .r(v1862ibus), .q(v1862obus), .dec(dec[1862]));
wire [data_w*2-1:0] v1863ibus;
wire [temp_w*2-1:0] v1863obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1863 (.l(l[1863*data_w +:data_w]), .r(v1863ibus), .q(v1863obus), .dec(dec[1863]));
wire [data_w*2-1:0] v1864ibus;
wire [temp_w*2-1:0] v1864obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1864 (.l(l[1864*data_w +:data_w]), .r(v1864ibus), .q(v1864obus), .dec(dec[1864]));
wire [data_w*2-1:0] v1865ibus;
wire [temp_w*2-1:0] v1865obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1865 (.l(l[1865*data_w +:data_w]), .r(v1865ibus), .q(v1865obus), .dec(dec[1865]));
wire [data_w*2-1:0] v1866ibus;
wire [temp_w*2-1:0] v1866obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1866 (.l(l[1866*data_w +:data_w]), .r(v1866ibus), .q(v1866obus), .dec(dec[1866]));
wire [data_w*2-1:0] v1867ibus;
wire [temp_w*2-1:0] v1867obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1867 (.l(l[1867*data_w +:data_w]), .r(v1867ibus), .q(v1867obus), .dec(dec[1867]));
wire [data_w*2-1:0] v1868ibus;
wire [temp_w*2-1:0] v1868obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1868 (.l(l[1868*data_w +:data_w]), .r(v1868ibus), .q(v1868obus), .dec(dec[1868]));
wire [data_w*2-1:0] v1869ibus;
wire [temp_w*2-1:0] v1869obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1869 (.l(l[1869*data_w +:data_w]), .r(v1869ibus), .q(v1869obus), .dec(dec[1869]));
wire [data_w*2-1:0] v1870ibus;
wire [temp_w*2-1:0] v1870obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1870 (.l(l[1870*data_w +:data_w]), .r(v1870ibus), .q(v1870obus), .dec(dec[1870]));
wire [data_w*2-1:0] v1871ibus;
wire [temp_w*2-1:0] v1871obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1871 (.l(l[1871*data_w +:data_w]), .r(v1871ibus), .q(v1871obus), .dec(dec[1871]));
wire [data_w*2-1:0] v1872ibus;
wire [temp_w*2-1:0] v1872obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1872 (.l(l[1872*data_w +:data_w]), .r(v1872ibus), .q(v1872obus), .dec(dec[1872]));
wire [data_w*2-1:0] v1873ibus;
wire [temp_w*2-1:0] v1873obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1873 (.l(l[1873*data_w +:data_w]), .r(v1873ibus), .q(v1873obus), .dec(dec[1873]));
wire [data_w*2-1:0] v1874ibus;
wire [temp_w*2-1:0] v1874obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1874 (.l(l[1874*data_w +:data_w]), .r(v1874ibus), .q(v1874obus), .dec(dec[1874]));
wire [data_w*2-1:0] v1875ibus;
wire [temp_w*2-1:0] v1875obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1875 (.l(l[1875*data_w +:data_w]), .r(v1875ibus), .q(v1875obus), .dec(dec[1875]));
wire [data_w*2-1:0] v1876ibus;
wire [temp_w*2-1:0] v1876obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1876 (.l(l[1876*data_w +:data_w]), .r(v1876ibus), .q(v1876obus), .dec(dec[1876]));
wire [data_w*2-1:0] v1877ibus;
wire [temp_w*2-1:0] v1877obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1877 (.l(l[1877*data_w +:data_w]), .r(v1877ibus), .q(v1877obus), .dec(dec[1877]));
wire [data_w*2-1:0] v1878ibus;
wire [temp_w*2-1:0] v1878obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1878 (.l(l[1878*data_w +:data_w]), .r(v1878ibus), .q(v1878obus), .dec(dec[1878]));
wire [data_w*2-1:0] v1879ibus;
wire [temp_w*2-1:0] v1879obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1879 (.l(l[1879*data_w +:data_w]), .r(v1879ibus), .q(v1879obus), .dec(dec[1879]));
wire [data_w*2-1:0] v1880ibus;
wire [temp_w*2-1:0] v1880obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1880 (.l(l[1880*data_w +:data_w]), .r(v1880ibus), .q(v1880obus), .dec(dec[1880]));
wire [data_w*2-1:0] v1881ibus;
wire [temp_w*2-1:0] v1881obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1881 (.l(l[1881*data_w +:data_w]), .r(v1881ibus), .q(v1881obus), .dec(dec[1881]));
wire [data_w*2-1:0] v1882ibus;
wire [temp_w*2-1:0] v1882obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1882 (.l(l[1882*data_w +:data_w]), .r(v1882ibus), .q(v1882obus), .dec(dec[1882]));
wire [data_w*2-1:0] v1883ibus;
wire [temp_w*2-1:0] v1883obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1883 (.l(l[1883*data_w +:data_w]), .r(v1883ibus), .q(v1883obus), .dec(dec[1883]));
wire [data_w*2-1:0] v1884ibus;
wire [temp_w*2-1:0] v1884obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1884 (.l(l[1884*data_w +:data_w]), .r(v1884ibus), .q(v1884obus), .dec(dec[1884]));
wire [data_w*2-1:0] v1885ibus;
wire [temp_w*2-1:0] v1885obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1885 (.l(l[1885*data_w +:data_w]), .r(v1885ibus), .q(v1885obus), .dec(dec[1885]));
wire [data_w*2-1:0] v1886ibus;
wire [temp_w*2-1:0] v1886obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1886 (.l(l[1886*data_w +:data_w]), .r(v1886ibus), .q(v1886obus), .dec(dec[1886]));
wire [data_w*2-1:0] v1887ibus;
wire [temp_w*2-1:0] v1887obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1887 (.l(l[1887*data_w +:data_w]), .r(v1887ibus), .q(v1887obus), .dec(dec[1887]));
wire [data_w*2-1:0] v1888ibus;
wire [temp_w*2-1:0] v1888obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1888 (.l(l[1888*data_w +:data_w]), .r(v1888ibus), .q(v1888obus), .dec(dec[1888]));
wire [data_w*2-1:0] v1889ibus;
wire [temp_w*2-1:0] v1889obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1889 (.l(l[1889*data_w +:data_w]), .r(v1889ibus), .q(v1889obus), .dec(dec[1889]));
wire [data_w*2-1:0] v1890ibus;
wire [temp_w*2-1:0] v1890obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1890 (.l(l[1890*data_w +:data_w]), .r(v1890ibus), .q(v1890obus), .dec(dec[1890]));
wire [data_w*2-1:0] v1891ibus;
wire [temp_w*2-1:0] v1891obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1891 (.l(l[1891*data_w +:data_w]), .r(v1891ibus), .q(v1891obus), .dec(dec[1891]));
wire [data_w*2-1:0] v1892ibus;
wire [temp_w*2-1:0] v1892obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1892 (.l(l[1892*data_w +:data_w]), .r(v1892ibus), .q(v1892obus), .dec(dec[1892]));
wire [data_w*2-1:0] v1893ibus;
wire [temp_w*2-1:0] v1893obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1893 (.l(l[1893*data_w +:data_w]), .r(v1893ibus), .q(v1893obus), .dec(dec[1893]));
wire [data_w*2-1:0] v1894ibus;
wire [temp_w*2-1:0] v1894obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1894 (.l(l[1894*data_w +:data_w]), .r(v1894ibus), .q(v1894obus), .dec(dec[1894]));
wire [data_w*2-1:0] v1895ibus;
wire [temp_w*2-1:0] v1895obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1895 (.l(l[1895*data_w +:data_w]), .r(v1895ibus), .q(v1895obus), .dec(dec[1895]));
wire [data_w*2-1:0] v1896ibus;
wire [temp_w*2-1:0] v1896obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1896 (.l(l[1896*data_w +:data_w]), .r(v1896ibus), .q(v1896obus), .dec(dec[1896]));
wire [data_w*2-1:0] v1897ibus;
wire [temp_w*2-1:0] v1897obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1897 (.l(l[1897*data_w +:data_w]), .r(v1897ibus), .q(v1897obus), .dec(dec[1897]));
wire [data_w*2-1:0] v1898ibus;
wire [temp_w*2-1:0] v1898obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1898 (.l(l[1898*data_w +:data_w]), .r(v1898ibus), .q(v1898obus), .dec(dec[1898]));
wire [data_w*2-1:0] v1899ibus;
wire [temp_w*2-1:0] v1899obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1899 (.l(l[1899*data_w +:data_w]), .r(v1899ibus), .q(v1899obus), .dec(dec[1899]));
wire [data_w*2-1:0] v1900ibus;
wire [temp_w*2-1:0] v1900obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1900 (.l(l[1900*data_w +:data_w]), .r(v1900ibus), .q(v1900obus), .dec(dec[1900]));
wire [data_w*2-1:0] v1901ibus;
wire [temp_w*2-1:0] v1901obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1901 (.l(l[1901*data_w +:data_w]), .r(v1901ibus), .q(v1901obus), .dec(dec[1901]));
wire [data_w*2-1:0] v1902ibus;
wire [temp_w*2-1:0] v1902obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1902 (.l(l[1902*data_w +:data_w]), .r(v1902ibus), .q(v1902obus), .dec(dec[1902]));
wire [data_w*2-1:0] v1903ibus;
wire [temp_w*2-1:0] v1903obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1903 (.l(l[1903*data_w +:data_w]), .r(v1903ibus), .q(v1903obus), .dec(dec[1903]));
wire [data_w*2-1:0] v1904ibus;
wire [temp_w*2-1:0] v1904obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1904 (.l(l[1904*data_w +:data_w]), .r(v1904ibus), .q(v1904obus), .dec(dec[1904]));
wire [data_w*2-1:0] v1905ibus;
wire [temp_w*2-1:0] v1905obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1905 (.l(l[1905*data_w +:data_w]), .r(v1905ibus), .q(v1905obus), .dec(dec[1905]));
wire [data_w*2-1:0] v1906ibus;
wire [temp_w*2-1:0] v1906obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1906 (.l(l[1906*data_w +:data_w]), .r(v1906ibus), .q(v1906obus), .dec(dec[1906]));
wire [data_w*2-1:0] v1907ibus;
wire [temp_w*2-1:0] v1907obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1907 (.l(l[1907*data_w +:data_w]), .r(v1907ibus), .q(v1907obus), .dec(dec[1907]));
wire [data_w*2-1:0] v1908ibus;
wire [temp_w*2-1:0] v1908obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1908 (.l(l[1908*data_w +:data_w]), .r(v1908ibus), .q(v1908obus), .dec(dec[1908]));
wire [data_w*2-1:0] v1909ibus;
wire [temp_w*2-1:0] v1909obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1909 (.l(l[1909*data_w +:data_w]), .r(v1909ibus), .q(v1909obus), .dec(dec[1909]));
wire [data_w*2-1:0] v1910ibus;
wire [temp_w*2-1:0] v1910obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1910 (.l(l[1910*data_w +:data_w]), .r(v1910ibus), .q(v1910obus), .dec(dec[1910]));
wire [data_w*2-1:0] v1911ibus;
wire [temp_w*2-1:0] v1911obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1911 (.l(l[1911*data_w +:data_w]), .r(v1911ibus), .q(v1911obus), .dec(dec[1911]));
wire [data_w*2-1:0] v1912ibus;
wire [temp_w*2-1:0] v1912obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1912 (.l(l[1912*data_w +:data_w]), .r(v1912ibus), .q(v1912obus), .dec(dec[1912]));
wire [data_w*2-1:0] v1913ibus;
wire [temp_w*2-1:0] v1913obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1913 (.l(l[1913*data_w +:data_w]), .r(v1913ibus), .q(v1913obus), .dec(dec[1913]));
wire [data_w*2-1:0] v1914ibus;
wire [temp_w*2-1:0] v1914obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1914 (.l(l[1914*data_w +:data_w]), .r(v1914ibus), .q(v1914obus), .dec(dec[1914]));
wire [data_w*2-1:0] v1915ibus;
wire [temp_w*2-1:0] v1915obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1915 (.l(l[1915*data_w +:data_w]), .r(v1915ibus), .q(v1915obus), .dec(dec[1915]));
wire [data_w*2-1:0] v1916ibus;
wire [temp_w*2-1:0] v1916obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1916 (.l(l[1916*data_w +:data_w]), .r(v1916ibus), .q(v1916obus), .dec(dec[1916]));
wire [data_w*2-1:0] v1917ibus;
wire [temp_w*2-1:0] v1917obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1917 (.l(l[1917*data_w +:data_w]), .r(v1917ibus), .q(v1917obus), .dec(dec[1917]));
wire [data_w*2-1:0] v1918ibus;
wire [temp_w*2-1:0] v1918obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1918 (.l(l[1918*data_w +:data_w]), .r(v1918ibus), .q(v1918obus), .dec(dec[1918]));
wire [data_w*2-1:0] v1919ibus;
wire [temp_w*2-1:0] v1919obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1919 (.l(l[1919*data_w +:data_w]), .r(v1919ibus), .q(v1919obus), .dec(dec[1919]));
wire [data_w*2-1:0] v1920ibus;
wire [temp_w*2-1:0] v1920obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1920 (.l(l[1920*data_w +:data_w]), .r(v1920ibus), .q(v1920obus), .dec(dec[1920]));
wire [data_w*2-1:0] v1921ibus;
wire [temp_w*2-1:0] v1921obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1921 (.l(l[1921*data_w +:data_w]), .r(v1921ibus), .q(v1921obus), .dec(dec[1921]));
wire [data_w*2-1:0] v1922ibus;
wire [temp_w*2-1:0] v1922obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1922 (.l(l[1922*data_w +:data_w]), .r(v1922ibus), .q(v1922obus), .dec(dec[1922]));
wire [data_w*2-1:0] v1923ibus;
wire [temp_w*2-1:0] v1923obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1923 (.l(l[1923*data_w +:data_w]), .r(v1923ibus), .q(v1923obus), .dec(dec[1923]));
wire [data_w*2-1:0] v1924ibus;
wire [temp_w*2-1:0] v1924obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1924 (.l(l[1924*data_w +:data_w]), .r(v1924ibus), .q(v1924obus), .dec(dec[1924]));
wire [data_w*2-1:0] v1925ibus;
wire [temp_w*2-1:0] v1925obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1925 (.l(l[1925*data_w +:data_w]), .r(v1925ibus), .q(v1925obus), .dec(dec[1925]));
wire [data_w*2-1:0] v1926ibus;
wire [temp_w*2-1:0] v1926obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1926 (.l(l[1926*data_w +:data_w]), .r(v1926ibus), .q(v1926obus), .dec(dec[1926]));
wire [data_w*2-1:0] v1927ibus;
wire [temp_w*2-1:0] v1927obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1927 (.l(l[1927*data_w +:data_w]), .r(v1927ibus), .q(v1927obus), .dec(dec[1927]));
wire [data_w*2-1:0] v1928ibus;
wire [temp_w*2-1:0] v1928obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1928 (.l(l[1928*data_w +:data_w]), .r(v1928ibus), .q(v1928obus), .dec(dec[1928]));
wire [data_w*2-1:0] v1929ibus;
wire [temp_w*2-1:0] v1929obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1929 (.l(l[1929*data_w +:data_w]), .r(v1929ibus), .q(v1929obus), .dec(dec[1929]));
wire [data_w*2-1:0] v1930ibus;
wire [temp_w*2-1:0] v1930obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1930 (.l(l[1930*data_w +:data_w]), .r(v1930ibus), .q(v1930obus), .dec(dec[1930]));
wire [data_w*2-1:0] v1931ibus;
wire [temp_w*2-1:0] v1931obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1931 (.l(l[1931*data_w +:data_w]), .r(v1931ibus), .q(v1931obus), .dec(dec[1931]));
wire [data_w*2-1:0] v1932ibus;
wire [temp_w*2-1:0] v1932obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1932 (.l(l[1932*data_w +:data_w]), .r(v1932ibus), .q(v1932obus), .dec(dec[1932]));
wire [data_w*2-1:0] v1933ibus;
wire [temp_w*2-1:0] v1933obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1933 (.l(l[1933*data_w +:data_w]), .r(v1933ibus), .q(v1933obus), .dec(dec[1933]));
wire [data_w*2-1:0] v1934ibus;
wire [temp_w*2-1:0] v1934obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1934 (.l(l[1934*data_w +:data_w]), .r(v1934ibus), .q(v1934obus), .dec(dec[1934]));
wire [data_w*2-1:0] v1935ibus;
wire [temp_w*2-1:0] v1935obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1935 (.l(l[1935*data_w +:data_w]), .r(v1935ibus), .q(v1935obus), .dec(dec[1935]));
wire [data_w*2-1:0] v1936ibus;
wire [temp_w*2-1:0] v1936obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1936 (.l(l[1936*data_w +:data_w]), .r(v1936ibus), .q(v1936obus), .dec(dec[1936]));
wire [data_w*2-1:0] v1937ibus;
wire [temp_w*2-1:0] v1937obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1937 (.l(l[1937*data_w +:data_w]), .r(v1937ibus), .q(v1937obus), .dec(dec[1937]));
wire [data_w*2-1:0] v1938ibus;
wire [temp_w*2-1:0] v1938obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1938 (.l(l[1938*data_w +:data_w]), .r(v1938ibus), .q(v1938obus), .dec(dec[1938]));
wire [data_w*2-1:0] v1939ibus;
wire [temp_w*2-1:0] v1939obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1939 (.l(l[1939*data_w +:data_w]), .r(v1939ibus), .q(v1939obus), .dec(dec[1939]));
wire [data_w*2-1:0] v1940ibus;
wire [temp_w*2-1:0] v1940obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1940 (.l(l[1940*data_w +:data_w]), .r(v1940ibus), .q(v1940obus), .dec(dec[1940]));
wire [data_w*2-1:0] v1941ibus;
wire [temp_w*2-1:0] v1941obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1941 (.l(l[1941*data_w +:data_w]), .r(v1941ibus), .q(v1941obus), .dec(dec[1941]));
wire [data_w*2-1:0] v1942ibus;
wire [temp_w*2-1:0] v1942obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1942 (.l(l[1942*data_w +:data_w]), .r(v1942ibus), .q(v1942obus), .dec(dec[1942]));
wire [data_w*2-1:0] v1943ibus;
wire [temp_w*2-1:0] v1943obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1943 (.l(l[1943*data_w +:data_w]), .r(v1943ibus), .q(v1943obus), .dec(dec[1943]));
wire [data_w*2-1:0] v1944ibus;
wire [temp_w*2-1:0] v1944obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1944 (.l(l[1944*data_w +:data_w]), .r(v1944ibus), .q(v1944obus), .dec(dec[1944]));
wire [data_w*2-1:0] v1945ibus;
wire [temp_w*2-1:0] v1945obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1945 (.l(l[1945*data_w +:data_w]), .r(v1945ibus), .q(v1945obus), .dec(dec[1945]));
wire [data_w*2-1:0] v1946ibus;
wire [temp_w*2-1:0] v1946obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1946 (.l(l[1946*data_w +:data_w]), .r(v1946ibus), .q(v1946obus), .dec(dec[1946]));
wire [data_w*2-1:0] v1947ibus;
wire [temp_w*2-1:0] v1947obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1947 (.l(l[1947*data_w +:data_w]), .r(v1947ibus), .q(v1947obus), .dec(dec[1947]));
wire [data_w*2-1:0] v1948ibus;
wire [temp_w*2-1:0] v1948obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1948 (.l(l[1948*data_w +:data_w]), .r(v1948ibus), .q(v1948obus), .dec(dec[1948]));
wire [data_w*2-1:0] v1949ibus;
wire [temp_w*2-1:0] v1949obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1949 (.l(l[1949*data_w +:data_w]), .r(v1949ibus), .q(v1949obus), .dec(dec[1949]));
wire [data_w*2-1:0] v1950ibus;
wire [temp_w*2-1:0] v1950obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1950 (.l(l[1950*data_w +:data_w]), .r(v1950ibus), .q(v1950obus), .dec(dec[1950]));
wire [data_w*2-1:0] v1951ibus;
wire [temp_w*2-1:0] v1951obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1951 (.l(l[1951*data_w +:data_w]), .r(v1951ibus), .q(v1951obus), .dec(dec[1951]));
wire [data_w*2-1:0] v1952ibus;
wire [temp_w*2-1:0] v1952obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1952 (.l(l[1952*data_w +:data_w]), .r(v1952ibus), .q(v1952obus), .dec(dec[1952]));
wire [data_w*2-1:0] v1953ibus;
wire [temp_w*2-1:0] v1953obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1953 (.l(l[1953*data_w +:data_w]), .r(v1953ibus), .q(v1953obus), .dec(dec[1953]));
wire [data_w*2-1:0] v1954ibus;
wire [temp_w*2-1:0] v1954obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1954 (.l(l[1954*data_w +:data_w]), .r(v1954ibus), .q(v1954obus), .dec(dec[1954]));
wire [data_w*2-1:0] v1955ibus;
wire [temp_w*2-1:0] v1955obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1955 (.l(l[1955*data_w +:data_w]), .r(v1955ibus), .q(v1955obus), .dec(dec[1955]));
wire [data_w*2-1:0] v1956ibus;
wire [temp_w*2-1:0] v1956obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1956 (.l(l[1956*data_w +:data_w]), .r(v1956ibus), .q(v1956obus), .dec(dec[1956]));
wire [data_w*2-1:0] v1957ibus;
wire [temp_w*2-1:0] v1957obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1957 (.l(l[1957*data_w +:data_w]), .r(v1957ibus), .q(v1957obus), .dec(dec[1957]));
wire [data_w*2-1:0] v1958ibus;
wire [temp_w*2-1:0] v1958obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1958 (.l(l[1958*data_w +:data_w]), .r(v1958ibus), .q(v1958obus), .dec(dec[1958]));
wire [data_w*2-1:0] v1959ibus;
wire [temp_w*2-1:0] v1959obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1959 (.l(l[1959*data_w +:data_w]), .r(v1959ibus), .q(v1959obus), .dec(dec[1959]));
wire [data_w*2-1:0] v1960ibus;
wire [temp_w*2-1:0] v1960obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1960 (.l(l[1960*data_w +:data_w]), .r(v1960ibus), .q(v1960obus), .dec(dec[1960]));
wire [data_w*2-1:0] v1961ibus;
wire [temp_w*2-1:0] v1961obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1961 (.l(l[1961*data_w +:data_w]), .r(v1961ibus), .q(v1961obus), .dec(dec[1961]));
wire [data_w*2-1:0] v1962ibus;
wire [temp_w*2-1:0] v1962obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1962 (.l(l[1962*data_w +:data_w]), .r(v1962ibus), .q(v1962obus), .dec(dec[1962]));
wire [data_w*2-1:0] v1963ibus;
wire [temp_w*2-1:0] v1963obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1963 (.l(l[1963*data_w +:data_w]), .r(v1963ibus), .q(v1963obus), .dec(dec[1963]));
wire [data_w*2-1:0] v1964ibus;
wire [temp_w*2-1:0] v1964obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1964 (.l(l[1964*data_w +:data_w]), .r(v1964ibus), .q(v1964obus), .dec(dec[1964]));
wire [data_w*2-1:0] v1965ibus;
wire [temp_w*2-1:0] v1965obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1965 (.l(l[1965*data_w +:data_w]), .r(v1965ibus), .q(v1965obus), .dec(dec[1965]));
wire [data_w*2-1:0] v1966ibus;
wire [temp_w*2-1:0] v1966obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1966 (.l(l[1966*data_w +:data_w]), .r(v1966ibus), .q(v1966obus), .dec(dec[1966]));
wire [data_w*2-1:0] v1967ibus;
wire [temp_w*2-1:0] v1967obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1967 (.l(l[1967*data_w +:data_w]), .r(v1967ibus), .q(v1967obus), .dec(dec[1967]));
wire [data_w*2-1:0] v1968ibus;
wire [temp_w*2-1:0] v1968obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1968 (.l(l[1968*data_w +:data_w]), .r(v1968ibus), .q(v1968obus), .dec(dec[1968]));
wire [data_w*2-1:0] v1969ibus;
wire [temp_w*2-1:0] v1969obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1969 (.l(l[1969*data_w +:data_w]), .r(v1969ibus), .q(v1969obus), .dec(dec[1969]));
wire [data_w*2-1:0] v1970ibus;
wire [temp_w*2-1:0] v1970obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1970 (.l(l[1970*data_w +:data_w]), .r(v1970ibus), .q(v1970obus), .dec(dec[1970]));
wire [data_w*2-1:0] v1971ibus;
wire [temp_w*2-1:0] v1971obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1971 (.l(l[1971*data_w +:data_w]), .r(v1971ibus), .q(v1971obus), .dec(dec[1971]));
wire [data_w*2-1:0] v1972ibus;
wire [temp_w*2-1:0] v1972obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1972 (.l(l[1972*data_w +:data_w]), .r(v1972ibus), .q(v1972obus), .dec(dec[1972]));
wire [data_w*2-1:0] v1973ibus;
wire [temp_w*2-1:0] v1973obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1973 (.l(l[1973*data_w +:data_w]), .r(v1973ibus), .q(v1973obus), .dec(dec[1973]));
wire [data_w*2-1:0] v1974ibus;
wire [temp_w*2-1:0] v1974obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1974 (.l(l[1974*data_w +:data_w]), .r(v1974ibus), .q(v1974obus), .dec(dec[1974]));
wire [data_w*2-1:0] v1975ibus;
wire [temp_w*2-1:0] v1975obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1975 (.l(l[1975*data_w +:data_w]), .r(v1975ibus), .q(v1975obus), .dec(dec[1975]));
wire [data_w*2-1:0] v1976ibus;
wire [temp_w*2-1:0] v1976obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1976 (.l(l[1976*data_w +:data_w]), .r(v1976ibus), .q(v1976obus), .dec(dec[1976]));
wire [data_w*2-1:0] v1977ibus;
wire [temp_w*2-1:0] v1977obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1977 (.l(l[1977*data_w +:data_w]), .r(v1977ibus), .q(v1977obus), .dec(dec[1977]));
wire [data_w*2-1:0] v1978ibus;
wire [temp_w*2-1:0] v1978obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1978 (.l(l[1978*data_w +:data_w]), .r(v1978ibus), .q(v1978obus), .dec(dec[1978]));
wire [data_w*2-1:0] v1979ibus;
wire [temp_w*2-1:0] v1979obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1979 (.l(l[1979*data_w +:data_w]), .r(v1979ibus), .q(v1979obus), .dec(dec[1979]));
wire [data_w*2-1:0] v1980ibus;
wire [temp_w*2-1:0] v1980obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1980 (.l(l[1980*data_w +:data_w]), .r(v1980ibus), .q(v1980obus), .dec(dec[1980]));
wire [data_w*2-1:0] v1981ibus;
wire [temp_w*2-1:0] v1981obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1981 (.l(l[1981*data_w +:data_w]), .r(v1981ibus), .q(v1981obus), .dec(dec[1981]));
wire [data_w*2-1:0] v1982ibus;
wire [temp_w*2-1:0] v1982obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1982 (.l(l[1982*data_w +:data_w]), .r(v1982ibus), .q(v1982obus), .dec(dec[1982]));
wire [data_w*2-1:0] v1983ibus;
wire [temp_w*2-1:0] v1983obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1983 (.l(l[1983*data_w +:data_w]), .r(v1983ibus), .q(v1983obus), .dec(dec[1983]));
wire [data_w*2-1:0] v1984ibus;
wire [temp_w*2-1:0] v1984obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1984 (.l(l[1984*data_w +:data_w]), .r(v1984ibus), .q(v1984obus), .dec(dec[1984]));
wire [data_w*2-1:0] v1985ibus;
wire [temp_w*2-1:0] v1985obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1985 (.l(l[1985*data_w +:data_w]), .r(v1985ibus), .q(v1985obus), .dec(dec[1985]));
wire [data_w*2-1:0] v1986ibus;
wire [temp_w*2-1:0] v1986obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1986 (.l(l[1986*data_w +:data_w]), .r(v1986ibus), .q(v1986obus), .dec(dec[1986]));
wire [data_w*2-1:0] v1987ibus;
wire [temp_w*2-1:0] v1987obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1987 (.l(l[1987*data_w +:data_w]), .r(v1987ibus), .q(v1987obus), .dec(dec[1987]));
wire [data_w*2-1:0] v1988ibus;
wire [temp_w*2-1:0] v1988obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1988 (.l(l[1988*data_w +:data_w]), .r(v1988ibus), .q(v1988obus), .dec(dec[1988]));
wire [data_w*2-1:0] v1989ibus;
wire [temp_w*2-1:0] v1989obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1989 (.l(l[1989*data_w +:data_w]), .r(v1989ibus), .q(v1989obus), .dec(dec[1989]));
wire [data_w*2-1:0] v1990ibus;
wire [temp_w*2-1:0] v1990obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1990 (.l(l[1990*data_w +:data_w]), .r(v1990ibus), .q(v1990obus), .dec(dec[1990]));
wire [data_w*2-1:0] v1991ibus;
wire [temp_w*2-1:0] v1991obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1991 (.l(l[1991*data_w +:data_w]), .r(v1991ibus), .q(v1991obus), .dec(dec[1991]));
wire [data_w*2-1:0] v1992ibus;
wire [temp_w*2-1:0] v1992obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1992 (.l(l[1992*data_w +:data_w]), .r(v1992ibus), .q(v1992obus), .dec(dec[1992]));
wire [data_w*2-1:0] v1993ibus;
wire [temp_w*2-1:0] v1993obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1993 (.l(l[1993*data_w +:data_w]), .r(v1993ibus), .q(v1993obus), .dec(dec[1993]));
wire [data_w*2-1:0] v1994ibus;
wire [temp_w*2-1:0] v1994obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1994 (.l(l[1994*data_w +:data_w]), .r(v1994ibus), .q(v1994obus), .dec(dec[1994]));
wire [data_w*2-1:0] v1995ibus;
wire [temp_w*2-1:0] v1995obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1995 (.l(l[1995*data_w +:data_w]), .r(v1995ibus), .q(v1995obus), .dec(dec[1995]));
wire [data_w*2-1:0] v1996ibus;
wire [temp_w*2-1:0] v1996obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1996 (.l(l[1996*data_w +:data_w]), .r(v1996ibus), .q(v1996obus), .dec(dec[1996]));
wire [data_w*2-1:0] v1997ibus;
wire [temp_w*2-1:0] v1997obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1997 (.l(l[1997*data_w +:data_w]), .r(v1997ibus), .q(v1997obus), .dec(dec[1997]));
wire [data_w*2-1:0] v1998ibus;
wire [temp_w*2-1:0] v1998obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1998 (.l(l[1998*data_w +:data_w]), .r(v1998ibus), .q(v1998obus), .dec(dec[1998]));
wire [data_w*2-1:0] v1999ibus;
wire [temp_w*2-1:0] v1999obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU1999 (.l(l[1999*data_w +:data_w]), .r(v1999ibus), .q(v1999obus), .dec(dec[1999]));
wire [data_w*2-1:0] v2000ibus;
wire [temp_w*2-1:0] v2000obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2000 (.l(l[2000*data_w +:data_w]), .r(v2000ibus), .q(v2000obus), .dec(dec[2000]));
wire [data_w*2-1:0] v2001ibus;
wire [temp_w*2-1:0] v2001obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2001 (.l(l[2001*data_w +:data_w]), .r(v2001ibus), .q(v2001obus), .dec(dec[2001]));
wire [data_w*2-1:0] v2002ibus;
wire [temp_w*2-1:0] v2002obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2002 (.l(l[2002*data_w +:data_w]), .r(v2002ibus), .q(v2002obus), .dec(dec[2002]));
wire [data_w*2-1:0] v2003ibus;
wire [temp_w*2-1:0] v2003obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2003 (.l(l[2003*data_w +:data_w]), .r(v2003ibus), .q(v2003obus), .dec(dec[2003]));
wire [data_w*2-1:0] v2004ibus;
wire [temp_w*2-1:0] v2004obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2004 (.l(l[2004*data_w +:data_w]), .r(v2004ibus), .q(v2004obus), .dec(dec[2004]));
wire [data_w*2-1:0] v2005ibus;
wire [temp_w*2-1:0] v2005obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2005 (.l(l[2005*data_w +:data_w]), .r(v2005ibus), .q(v2005obus), .dec(dec[2005]));
wire [data_w*2-1:0] v2006ibus;
wire [temp_w*2-1:0] v2006obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2006 (.l(l[2006*data_w +:data_w]), .r(v2006ibus), .q(v2006obus), .dec(dec[2006]));
wire [data_w*2-1:0] v2007ibus;
wire [temp_w*2-1:0] v2007obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2007 (.l(l[2007*data_w +:data_w]), .r(v2007ibus), .q(v2007obus), .dec(dec[2007]));
wire [data_w*2-1:0] v2008ibus;
wire [temp_w*2-1:0] v2008obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2008 (.l(l[2008*data_w +:data_w]), .r(v2008ibus), .q(v2008obus), .dec(dec[2008]));
wire [data_w*2-1:0] v2009ibus;
wire [temp_w*2-1:0] v2009obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2009 (.l(l[2009*data_w +:data_w]), .r(v2009ibus), .q(v2009obus), .dec(dec[2009]));
wire [data_w*2-1:0] v2010ibus;
wire [temp_w*2-1:0] v2010obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2010 (.l(l[2010*data_w +:data_w]), .r(v2010ibus), .q(v2010obus), .dec(dec[2010]));
wire [data_w*2-1:0] v2011ibus;
wire [temp_w*2-1:0] v2011obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2011 (.l(l[2011*data_w +:data_w]), .r(v2011ibus), .q(v2011obus), .dec(dec[2011]));
wire [data_w*2-1:0] v2012ibus;
wire [temp_w*2-1:0] v2012obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2012 (.l(l[2012*data_w +:data_w]), .r(v2012ibus), .q(v2012obus), .dec(dec[2012]));
wire [data_w*2-1:0] v2013ibus;
wire [temp_w*2-1:0] v2013obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2013 (.l(l[2013*data_w +:data_w]), .r(v2013ibus), .q(v2013obus), .dec(dec[2013]));
wire [data_w*2-1:0] v2014ibus;
wire [temp_w*2-1:0] v2014obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2014 (.l(l[2014*data_w +:data_w]), .r(v2014ibus), .q(v2014obus), .dec(dec[2014]));
wire [data_w*2-1:0] v2015ibus;
wire [temp_w*2-1:0] v2015obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2015 (.l(l[2015*data_w +:data_w]), .r(v2015ibus), .q(v2015obus), .dec(dec[2015]));
wire [data_w*2-1:0] v2016ibus;
wire [temp_w*2-1:0] v2016obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2016 (.l(l[2016*data_w +:data_w]), .r(v2016ibus), .q(v2016obus), .dec(dec[2016]));
wire [data_w*2-1:0] v2017ibus;
wire [temp_w*2-1:0] v2017obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2017 (.l(l[2017*data_w +:data_w]), .r(v2017ibus), .q(v2017obus), .dec(dec[2017]));
wire [data_w*2-1:0] v2018ibus;
wire [temp_w*2-1:0] v2018obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2018 (.l(l[2018*data_w +:data_w]), .r(v2018ibus), .q(v2018obus), .dec(dec[2018]));
wire [data_w*2-1:0] v2019ibus;
wire [temp_w*2-1:0] v2019obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2019 (.l(l[2019*data_w +:data_w]), .r(v2019ibus), .q(v2019obus), .dec(dec[2019]));
wire [data_w*2-1:0] v2020ibus;
wire [temp_w*2-1:0] v2020obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2020 (.l(l[2020*data_w +:data_w]), .r(v2020ibus), .q(v2020obus), .dec(dec[2020]));
wire [data_w*2-1:0] v2021ibus;
wire [temp_w*2-1:0] v2021obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2021 (.l(l[2021*data_w +:data_w]), .r(v2021ibus), .q(v2021obus), .dec(dec[2021]));
wire [data_w*2-1:0] v2022ibus;
wire [temp_w*2-1:0] v2022obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2022 (.l(l[2022*data_w +:data_w]), .r(v2022ibus), .q(v2022obus), .dec(dec[2022]));
wire [data_w*2-1:0] v2023ibus;
wire [temp_w*2-1:0] v2023obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2023 (.l(l[2023*data_w +:data_w]), .r(v2023ibus), .q(v2023obus), .dec(dec[2023]));
wire [data_w*2-1:0] v2024ibus;
wire [temp_w*2-1:0] v2024obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2024 (.l(l[2024*data_w +:data_w]), .r(v2024ibus), .q(v2024obus), .dec(dec[2024]));
wire [data_w*2-1:0] v2025ibus;
wire [temp_w*2-1:0] v2025obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2025 (.l(l[2025*data_w +:data_w]), .r(v2025ibus), .q(v2025obus), .dec(dec[2025]));
wire [data_w*2-1:0] v2026ibus;
wire [temp_w*2-1:0] v2026obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2026 (.l(l[2026*data_w +:data_w]), .r(v2026ibus), .q(v2026obus), .dec(dec[2026]));
wire [data_w*2-1:0] v2027ibus;
wire [temp_w*2-1:0] v2027obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2027 (.l(l[2027*data_w +:data_w]), .r(v2027ibus), .q(v2027obus), .dec(dec[2027]));
wire [data_w*2-1:0] v2028ibus;
wire [temp_w*2-1:0] v2028obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2028 (.l(l[2028*data_w +:data_w]), .r(v2028ibus), .q(v2028obus), .dec(dec[2028]));
wire [data_w*2-1:0] v2029ibus;
wire [temp_w*2-1:0] v2029obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2029 (.l(l[2029*data_w +:data_w]), .r(v2029ibus), .q(v2029obus), .dec(dec[2029]));
wire [data_w*2-1:0] v2030ibus;
wire [temp_w*2-1:0] v2030obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2030 (.l(l[2030*data_w +:data_w]), .r(v2030ibus), .q(v2030obus), .dec(dec[2030]));
wire [data_w*2-1:0] v2031ibus;
wire [temp_w*2-1:0] v2031obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2031 (.l(l[2031*data_w +:data_w]), .r(v2031ibus), .q(v2031obus), .dec(dec[2031]));
wire [data_w*2-1:0] v2032ibus;
wire [temp_w*2-1:0] v2032obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2032 (.l(l[2032*data_w +:data_w]), .r(v2032ibus), .q(v2032obus), .dec(dec[2032]));
wire [data_w*2-1:0] v2033ibus;
wire [temp_w*2-1:0] v2033obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2033 (.l(l[2033*data_w +:data_w]), .r(v2033ibus), .q(v2033obus), .dec(dec[2033]));
wire [data_w*2-1:0] v2034ibus;
wire [temp_w*2-1:0] v2034obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2034 (.l(l[2034*data_w +:data_w]), .r(v2034ibus), .q(v2034obus), .dec(dec[2034]));
wire [data_w*2-1:0] v2035ibus;
wire [temp_w*2-1:0] v2035obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2035 (.l(l[2035*data_w +:data_w]), .r(v2035ibus), .q(v2035obus), .dec(dec[2035]));
wire [data_w*2-1:0] v2036ibus;
wire [temp_w*2-1:0] v2036obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2036 (.l(l[2036*data_w +:data_w]), .r(v2036ibus), .q(v2036obus), .dec(dec[2036]));
wire [data_w*2-1:0] v2037ibus;
wire [temp_w*2-1:0] v2037obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2037 (.l(l[2037*data_w +:data_w]), .r(v2037ibus), .q(v2037obus), .dec(dec[2037]));
wire [data_w*2-1:0] v2038ibus;
wire [temp_w*2-1:0] v2038obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2038 (.l(l[2038*data_w +:data_w]), .r(v2038ibus), .q(v2038obus), .dec(dec[2038]));
wire [data_w*2-1:0] v2039ibus;
wire [temp_w*2-1:0] v2039obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2039 (.l(l[2039*data_w +:data_w]), .r(v2039ibus), .q(v2039obus), .dec(dec[2039]));
wire [data_w*2-1:0] v2040ibus;
wire [temp_w*2-1:0] v2040obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2040 (.l(l[2040*data_w +:data_w]), .r(v2040ibus), .q(v2040obus), .dec(dec[2040]));
wire [data_w*2-1:0] v2041ibus;
wire [temp_w*2-1:0] v2041obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2041 (.l(l[2041*data_w +:data_w]), .r(v2041ibus), .q(v2041obus), .dec(dec[2041]));
wire [data_w*2-1:0] v2042ibus;
wire [temp_w*2-1:0] v2042obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2042 (.l(l[2042*data_w +:data_w]), .r(v2042ibus), .q(v2042obus), .dec(dec[2042]));
wire [data_w*2-1:0] v2043ibus;
wire [temp_w*2-1:0] v2043obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2043 (.l(l[2043*data_w +:data_w]), .r(v2043ibus), .q(v2043obus), .dec(dec[2043]));
wire [data_w*2-1:0] v2044ibus;
wire [temp_w*2-1:0] v2044obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2044 (.l(l[2044*data_w +:data_w]), .r(v2044ibus), .q(v2044obus), .dec(dec[2044]));
wire [data_w*2-1:0] v2045ibus;
wire [temp_w*2-1:0] v2045obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2045 (.l(l[2045*data_w +:data_w]), .r(v2045ibus), .q(v2045obus), .dec(dec[2045]));
wire [data_w*2-1:0] v2046ibus;
wire [temp_w*2-1:0] v2046obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2046 (.l(l[2046*data_w +:data_w]), .r(v2046ibus), .q(v2046obus), .dec(dec[2046]));
wire [data_w*2-1:0] v2047ibus;
wire [temp_w*2-1:0] v2047obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2047 (.l(l[2047*data_w +:data_w]), .r(v2047ibus), .q(v2047obus), .dec(dec[2047]));
wire [data_w*2-1:0] v2048ibus;
wire [temp_w*2-1:0] v2048obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2048 (.l(l[2048*data_w +:data_w]), .r(v2048ibus), .q(v2048obus), .dec(dec[2048]));
wire [data_w*2-1:0] v2049ibus;
wire [temp_w*2-1:0] v2049obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2049 (.l(l[2049*data_w +:data_w]), .r(v2049ibus), .q(v2049obus), .dec(dec[2049]));
wire [data_w*2-1:0] v2050ibus;
wire [temp_w*2-1:0] v2050obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2050 (.l(l[2050*data_w +:data_w]), .r(v2050ibus), .q(v2050obus), .dec(dec[2050]));
wire [data_w*2-1:0] v2051ibus;
wire [temp_w*2-1:0] v2051obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2051 (.l(l[2051*data_w +:data_w]), .r(v2051ibus), .q(v2051obus), .dec(dec[2051]));
wire [data_w*2-1:0] v2052ibus;
wire [temp_w*2-1:0] v2052obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2052 (.l(l[2052*data_w +:data_w]), .r(v2052ibus), .q(v2052obus), .dec(dec[2052]));
wire [data_w*2-1:0] v2053ibus;
wire [temp_w*2-1:0] v2053obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2053 (.l(l[2053*data_w +:data_w]), .r(v2053ibus), .q(v2053obus), .dec(dec[2053]));
wire [data_w*2-1:0] v2054ibus;
wire [temp_w*2-1:0] v2054obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2054 (.l(l[2054*data_w +:data_w]), .r(v2054ibus), .q(v2054obus), .dec(dec[2054]));
wire [data_w*2-1:0] v2055ibus;
wire [temp_w*2-1:0] v2055obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2055 (.l(l[2055*data_w +:data_w]), .r(v2055ibus), .q(v2055obus), .dec(dec[2055]));
wire [data_w*2-1:0] v2056ibus;
wire [temp_w*2-1:0] v2056obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2056 (.l(l[2056*data_w +:data_w]), .r(v2056ibus), .q(v2056obus), .dec(dec[2056]));
wire [data_w*2-1:0] v2057ibus;
wire [temp_w*2-1:0] v2057obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2057 (.l(l[2057*data_w +:data_w]), .r(v2057ibus), .q(v2057obus), .dec(dec[2057]));
wire [data_w*2-1:0] v2058ibus;
wire [temp_w*2-1:0] v2058obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2058 (.l(l[2058*data_w +:data_w]), .r(v2058ibus), .q(v2058obus), .dec(dec[2058]));
wire [data_w*2-1:0] v2059ibus;
wire [temp_w*2-1:0] v2059obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2059 (.l(l[2059*data_w +:data_w]), .r(v2059ibus), .q(v2059obus), .dec(dec[2059]));
wire [data_w*2-1:0] v2060ibus;
wire [temp_w*2-1:0] v2060obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2060 (.l(l[2060*data_w +:data_w]), .r(v2060ibus), .q(v2060obus), .dec(dec[2060]));
wire [data_w*2-1:0] v2061ibus;
wire [temp_w*2-1:0] v2061obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2061 (.l(l[2061*data_w +:data_w]), .r(v2061ibus), .q(v2061obus), .dec(dec[2061]));
wire [data_w*2-1:0] v2062ibus;
wire [temp_w*2-1:0] v2062obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2062 (.l(l[2062*data_w +:data_w]), .r(v2062ibus), .q(v2062obus), .dec(dec[2062]));
wire [data_w*2-1:0] v2063ibus;
wire [temp_w*2-1:0] v2063obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2063 (.l(l[2063*data_w +:data_w]), .r(v2063ibus), .q(v2063obus), .dec(dec[2063]));
wire [data_w*2-1:0] v2064ibus;
wire [temp_w*2-1:0] v2064obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2064 (.l(l[2064*data_w +:data_w]), .r(v2064ibus), .q(v2064obus), .dec(dec[2064]));
wire [data_w*2-1:0] v2065ibus;
wire [temp_w*2-1:0] v2065obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2065 (.l(l[2065*data_w +:data_w]), .r(v2065ibus), .q(v2065obus), .dec(dec[2065]));
wire [data_w*2-1:0] v2066ibus;
wire [temp_w*2-1:0] v2066obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2066 (.l(l[2066*data_w +:data_w]), .r(v2066ibus), .q(v2066obus), .dec(dec[2066]));
wire [data_w*2-1:0] v2067ibus;
wire [temp_w*2-1:0] v2067obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2067 (.l(l[2067*data_w +:data_w]), .r(v2067ibus), .q(v2067obus), .dec(dec[2067]));
wire [data_w*2-1:0] v2068ibus;
wire [temp_w*2-1:0] v2068obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2068 (.l(l[2068*data_w +:data_w]), .r(v2068ibus), .q(v2068obus), .dec(dec[2068]));
wire [data_w*2-1:0] v2069ibus;
wire [temp_w*2-1:0] v2069obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2069 (.l(l[2069*data_w +:data_w]), .r(v2069ibus), .q(v2069obus), .dec(dec[2069]));
wire [data_w*2-1:0] v2070ibus;
wire [temp_w*2-1:0] v2070obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2070 (.l(l[2070*data_w +:data_w]), .r(v2070ibus), .q(v2070obus), .dec(dec[2070]));
wire [data_w*2-1:0] v2071ibus;
wire [temp_w*2-1:0] v2071obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2071 (.l(l[2071*data_w +:data_w]), .r(v2071ibus), .q(v2071obus), .dec(dec[2071]));
wire [data_w*2-1:0] v2072ibus;
wire [temp_w*2-1:0] v2072obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2072 (.l(l[2072*data_w +:data_w]), .r(v2072ibus), .q(v2072obus), .dec(dec[2072]));
wire [data_w*2-1:0] v2073ibus;
wire [temp_w*2-1:0] v2073obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2073 (.l(l[2073*data_w +:data_w]), .r(v2073ibus), .q(v2073obus), .dec(dec[2073]));
wire [data_w*2-1:0] v2074ibus;
wire [temp_w*2-1:0] v2074obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2074 (.l(l[2074*data_w +:data_w]), .r(v2074ibus), .q(v2074obus), .dec(dec[2074]));
wire [data_w*2-1:0] v2075ibus;
wire [temp_w*2-1:0] v2075obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2075 (.l(l[2075*data_w +:data_w]), .r(v2075ibus), .q(v2075obus), .dec(dec[2075]));
wire [data_w*2-1:0] v2076ibus;
wire [temp_w*2-1:0] v2076obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2076 (.l(l[2076*data_w +:data_w]), .r(v2076ibus), .q(v2076obus), .dec(dec[2076]));
wire [data_w*2-1:0] v2077ibus;
wire [temp_w*2-1:0] v2077obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2077 (.l(l[2077*data_w +:data_w]), .r(v2077ibus), .q(v2077obus), .dec(dec[2077]));
wire [data_w*2-1:0] v2078ibus;
wire [temp_w*2-1:0] v2078obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2078 (.l(l[2078*data_w +:data_w]), .r(v2078ibus), .q(v2078obus), .dec(dec[2078]));
wire [data_w*2-1:0] v2079ibus;
wire [temp_w*2-1:0] v2079obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2079 (.l(l[2079*data_w +:data_w]), .r(v2079ibus), .q(v2079obus), .dec(dec[2079]));
wire [data_w*2-1:0] v2080ibus;
wire [temp_w*2-1:0] v2080obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2080 (.l(l[2080*data_w +:data_w]), .r(v2080ibus), .q(v2080obus), .dec(dec[2080]));
wire [data_w*2-1:0] v2081ibus;
wire [temp_w*2-1:0] v2081obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2081 (.l(l[2081*data_w +:data_w]), .r(v2081ibus), .q(v2081obus), .dec(dec[2081]));
wire [data_w*2-1:0] v2082ibus;
wire [temp_w*2-1:0] v2082obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2082 (.l(l[2082*data_w +:data_w]), .r(v2082ibus), .q(v2082obus), .dec(dec[2082]));
wire [data_w*2-1:0] v2083ibus;
wire [temp_w*2-1:0] v2083obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2083 (.l(l[2083*data_w +:data_w]), .r(v2083ibus), .q(v2083obus), .dec(dec[2083]));
wire [data_w*2-1:0] v2084ibus;
wire [temp_w*2-1:0] v2084obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2084 (.l(l[2084*data_w +:data_w]), .r(v2084ibus), .q(v2084obus), .dec(dec[2084]));
wire [data_w*2-1:0] v2085ibus;
wire [temp_w*2-1:0] v2085obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2085 (.l(l[2085*data_w +:data_w]), .r(v2085ibus), .q(v2085obus), .dec(dec[2085]));
wire [data_w*2-1:0] v2086ibus;
wire [temp_w*2-1:0] v2086obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2086 (.l(l[2086*data_w +:data_w]), .r(v2086ibus), .q(v2086obus), .dec(dec[2086]));
wire [data_w*2-1:0] v2087ibus;
wire [temp_w*2-1:0] v2087obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2087 (.l(l[2087*data_w +:data_w]), .r(v2087ibus), .q(v2087obus), .dec(dec[2087]));
wire [data_w*2-1:0] v2088ibus;
wire [temp_w*2-1:0] v2088obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2088 (.l(l[2088*data_w +:data_w]), .r(v2088ibus), .q(v2088obus), .dec(dec[2088]));
wire [data_w*2-1:0] v2089ibus;
wire [temp_w*2-1:0] v2089obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2089 (.l(l[2089*data_w +:data_w]), .r(v2089ibus), .q(v2089obus), .dec(dec[2089]));
wire [data_w*2-1:0] v2090ibus;
wire [temp_w*2-1:0] v2090obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2090 (.l(l[2090*data_w +:data_w]), .r(v2090ibus), .q(v2090obus), .dec(dec[2090]));
wire [data_w*2-1:0] v2091ibus;
wire [temp_w*2-1:0] v2091obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2091 (.l(l[2091*data_w +:data_w]), .r(v2091ibus), .q(v2091obus), .dec(dec[2091]));
wire [data_w*2-1:0] v2092ibus;
wire [temp_w*2-1:0] v2092obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2092 (.l(l[2092*data_w +:data_w]), .r(v2092ibus), .q(v2092obus), .dec(dec[2092]));
wire [data_w*2-1:0] v2093ibus;
wire [temp_w*2-1:0] v2093obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2093 (.l(l[2093*data_w +:data_w]), .r(v2093ibus), .q(v2093obus), .dec(dec[2093]));
wire [data_w*2-1:0] v2094ibus;
wire [temp_w*2-1:0] v2094obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2094 (.l(l[2094*data_w +:data_w]), .r(v2094ibus), .q(v2094obus), .dec(dec[2094]));
wire [data_w*2-1:0] v2095ibus;
wire [temp_w*2-1:0] v2095obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2095 (.l(l[2095*data_w +:data_w]), .r(v2095ibus), .q(v2095obus), .dec(dec[2095]));
wire [data_w*2-1:0] v2096ibus;
wire [temp_w*2-1:0] v2096obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2096 (.l(l[2096*data_w +:data_w]), .r(v2096ibus), .q(v2096obus), .dec(dec[2096]));
wire [data_w*2-1:0] v2097ibus;
wire [temp_w*2-1:0] v2097obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2097 (.l(l[2097*data_w +:data_w]), .r(v2097ibus), .q(v2097obus), .dec(dec[2097]));
wire [data_w*2-1:0] v2098ibus;
wire [temp_w*2-1:0] v2098obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2098 (.l(l[2098*data_w +:data_w]), .r(v2098ibus), .q(v2098obus), .dec(dec[2098]));
wire [data_w*2-1:0] v2099ibus;
wire [temp_w*2-1:0] v2099obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2099 (.l(l[2099*data_w +:data_w]), .r(v2099ibus), .q(v2099obus), .dec(dec[2099]));
wire [data_w*2-1:0] v2100ibus;
wire [temp_w*2-1:0] v2100obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2100 (.l(l[2100*data_w +:data_w]), .r(v2100ibus), .q(v2100obus), .dec(dec[2100]));
wire [data_w*2-1:0] v2101ibus;
wire [temp_w*2-1:0] v2101obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2101 (.l(l[2101*data_w +:data_w]), .r(v2101ibus), .q(v2101obus), .dec(dec[2101]));
wire [data_w*2-1:0] v2102ibus;
wire [temp_w*2-1:0] v2102obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2102 (.l(l[2102*data_w +:data_w]), .r(v2102ibus), .q(v2102obus), .dec(dec[2102]));
wire [data_w*2-1:0] v2103ibus;
wire [temp_w*2-1:0] v2103obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2103 (.l(l[2103*data_w +:data_w]), .r(v2103ibus), .q(v2103obus), .dec(dec[2103]));
wire [data_w*2-1:0] v2104ibus;
wire [temp_w*2-1:0] v2104obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2104 (.l(l[2104*data_w +:data_w]), .r(v2104ibus), .q(v2104obus), .dec(dec[2104]));
wire [data_w*2-1:0] v2105ibus;
wire [temp_w*2-1:0] v2105obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2105 (.l(l[2105*data_w +:data_w]), .r(v2105ibus), .q(v2105obus), .dec(dec[2105]));
wire [data_w*2-1:0] v2106ibus;
wire [temp_w*2-1:0] v2106obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2106 (.l(l[2106*data_w +:data_w]), .r(v2106ibus), .q(v2106obus), .dec(dec[2106]));
wire [data_w*2-1:0] v2107ibus;
wire [temp_w*2-1:0] v2107obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2107 (.l(l[2107*data_w +:data_w]), .r(v2107ibus), .q(v2107obus), .dec(dec[2107]));
wire [data_w*2-1:0] v2108ibus;
wire [temp_w*2-1:0] v2108obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2108 (.l(l[2108*data_w +:data_w]), .r(v2108ibus), .q(v2108obus), .dec(dec[2108]));
wire [data_w*2-1:0] v2109ibus;
wire [temp_w*2-1:0] v2109obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2109 (.l(l[2109*data_w +:data_w]), .r(v2109ibus), .q(v2109obus), .dec(dec[2109]));
wire [data_w*2-1:0] v2110ibus;
wire [temp_w*2-1:0] v2110obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2110 (.l(l[2110*data_w +:data_w]), .r(v2110ibus), .q(v2110obus), .dec(dec[2110]));
wire [data_w*2-1:0] v2111ibus;
wire [temp_w*2-1:0] v2111obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2111 (.l(l[2111*data_w +:data_w]), .r(v2111ibus), .q(v2111obus), .dec(dec[2111]));
wire [data_w*2-1:0] v2112ibus;
wire [temp_w*2-1:0] v2112obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2112 (.l(l[2112*data_w +:data_w]), .r(v2112ibus), .q(v2112obus), .dec(dec[2112]));
wire [data_w*2-1:0] v2113ibus;
wire [temp_w*2-1:0] v2113obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2113 (.l(l[2113*data_w +:data_w]), .r(v2113ibus), .q(v2113obus), .dec(dec[2113]));
wire [data_w*2-1:0] v2114ibus;
wire [temp_w*2-1:0] v2114obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2114 (.l(l[2114*data_w +:data_w]), .r(v2114ibus), .q(v2114obus), .dec(dec[2114]));
wire [data_w*2-1:0] v2115ibus;
wire [temp_w*2-1:0] v2115obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2115 (.l(l[2115*data_w +:data_w]), .r(v2115ibus), .q(v2115obus), .dec(dec[2115]));
wire [data_w*2-1:0] v2116ibus;
wire [temp_w*2-1:0] v2116obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2116 (.l(l[2116*data_w +:data_w]), .r(v2116ibus), .q(v2116obus), .dec(dec[2116]));
wire [data_w*2-1:0] v2117ibus;
wire [temp_w*2-1:0] v2117obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2117 (.l(l[2117*data_w +:data_w]), .r(v2117ibus), .q(v2117obus), .dec(dec[2117]));
wire [data_w*2-1:0] v2118ibus;
wire [temp_w*2-1:0] v2118obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2118 (.l(l[2118*data_w +:data_w]), .r(v2118ibus), .q(v2118obus), .dec(dec[2118]));
wire [data_w*2-1:0] v2119ibus;
wire [temp_w*2-1:0] v2119obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2119 (.l(l[2119*data_w +:data_w]), .r(v2119ibus), .q(v2119obus), .dec(dec[2119]));
wire [data_w*2-1:0] v2120ibus;
wire [temp_w*2-1:0] v2120obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2120 (.l(l[2120*data_w +:data_w]), .r(v2120ibus), .q(v2120obus), .dec(dec[2120]));
wire [data_w*2-1:0] v2121ibus;
wire [temp_w*2-1:0] v2121obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2121 (.l(l[2121*data_w +:data_w]), .r(v2121ibus), .q(v2121obus), .dec(dec[2121]));
wire [data_w*2-1:0] v2122ibus;
wire [temp_w*2-1:0] v2122obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2122 (.l(l[2122*data_w +:data_w]), .r(v2122ibus), .q(v2122obus), .dec(dec[2122]));
wire [data_w*2-1:0] v2123ibus;
wire [temp_w*2-1:0] v2123obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2123 (.l(l[2123*data_w +:data_w]), .r(v2123ibus), .q(v2123obus), .dec(dec[2123]));
wire [data_w*2-1:0] v2124ibus;
wire [temp_w*2-1:0] v2124obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2124 (.l(l[2124*data_w +:data_w]), .r(v2124ibus), .q(v2124obus), .dec(dec[2124]));
wire [data_w*2-1:0] v2125ibus;
wire [temp_w*2-1:0] v2125obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2125 (.l(l[2125*data_w +:data_w]), .r(v2125ibus), .q(v2125obus), .dec(dec[2125]));
wire [data_w*2-1:0] v2126ibus;
wire [temp_w*2-1:0] v2126obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2126 (.l(l[2126*data_w +:data_w]), .r(v2126ibus), .q(v2126obus), .dec(dec[2126]));
wire [data_w*2-1:0] v2127ibus;
wire [temp_w*2-1:0] v2127obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2127 (.l(l[2127*data_w +:data_w]), .r(v2127ibus), .q(v2127obus), .dec(dec[2127]));
wire [data_w*2-1:0] v2128ibus;
wire [temp_w*2-1:0] v2128obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2128 (.l(l[2128*data_w +:data_w]), .r(v2128ibus), .q(v2128obus), .dec(dec[2128]));
wire [data_w*2-1:0] v2129ibus;
wire [temp_w*2-1:0] v2129obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2129 (.l(l[2129*data_w +:data_w]), .r(v2129ibus), .q(v2129obus), .dec(dec[2129]));
wire [data_w*2-1:0] v2130ibus;
wire [temp_w*2-1:0] v2130obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2130 (.l(l[2130*data_w +:data_w]), .r(v2130ibus), .q(v2130obus), .dec(dec[2130]));
wire [data_w*2-1:0] v2131ibus;
wire [temp_w*2-1:0] v2131obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2131 (.l(l[2131*data_w +:data_w]), .r(v2131ibus), .q(v2131obus), .dec(dec[2131]));
wire [data_w*2-1:0] v2132ibus;
wire [temp_w*2-1:0] v2132obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2132 (.l(l[2132*data_w +:data_w]), .r(v2132ibus), .q(v2132obus), .dec(dec[2132]));
wire [data_w*2-1:0] v2133ibus;
wire [temp_w*2-1:0] v2133obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2133 (.l(l[2133*data_w +:data_w]), .r(v2133ibus), .q(v2133obus), .dec(dec[2133]));
wire [data_w*2-1:0] v2134ibus;
wire [temp_w*2-1:0] v2134obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2134 (.l(l[2134*data_w +:data_w]), .r(v2134ibus), .q(v2134obus), .dec(dec[2134]));
wire [data_w*2-1:0] v2135ibus;
wire [temp_w*2-1:0] v2135obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2135 (.l(l[2135*data_w +:data_w]), .r(v2135ibus), .q(v2135obus), .dec(dec[2135]));
wire [data_w*2-1:0] v2136ibus;
wire [temp_w*2-1:0] v2136obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2136 (.l(l[2136*data_w +:data_w]), .r(v2136ibus), .q(v2136obus), .dec(dec[2136]));
wire [data_w*2-1:0] v2137ibus;
wire [temp_w*2-1:0] v2137obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2137 (.l(l[2137*data_w +:data_w]), .r(v2137ibus), .q(v2137obus), .dec(dec[2137]));
wire [data_w*2-1:0] v2138ibus;
wire [temp_w*2-1:0] v2138obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2138 (.l(l[2138*data_w +:data_w]), .r(v2138ibus), .q(v2138obus), .dec(dec[2138]));
wire [data_w*2-1:0] v2139ibus;
wire [temp_w*2-1:0] v2139obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2139 (.l(l[2139*data_w +:data_w]), .r(v2139ibus), .q(v2139obus), .dec(dec[2139]));
wire [data_w*2-1:0] v2140ibus;
wire [temp_w*2-1:0] v2140obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2140 (.l(l[2140*data_w +:data_w]), .r(v2140ibus), .q(v2140obus), .dec(dec[2140]));
wire [data_w*2-1:0] v2141ibus;
wire [temp_w*2-1:0] v2141obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2141 (.l(l[2141*data_w +:data_w]), .r(v2141ibus), .q(v2141obus), .dec(dec[2141]));
wire [data_w*2-1:0] v2142ibus;
wire [temp_w*2-1:0] v2142obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2142 (.l(l[2142*data_w +:data_w]), .r(v2142ibus), .q(v2142obus), .dec(dec[2142]));
wire [data_w*2-1:0] v2143ibus;
wire [temp_w*2-1:0] v2143obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2143 (.l(l[2143*data_w +:data_w]), .r(v2143ibus), .q(v2143obus), .dec(dec[2143]));
wire [data_w*2-1:0] v2144ibus;
wire [temp_w*2-1:0] v2144obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2144 (.l(l[2144*data_w +:data_w]), .r(v2144ibus), .q(v2144obus), .dec(dec[2144]));
wire [data_w*2-1:0] v2145ibus;
wire [temp_w*2-1:0] v2145obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2145 (.l(l[2145*data_w +:data_w]), .r(v2145ibus), .q(v2145obus), .dec(dec[2145]));
wire [data_w*2-1:0] v2146ibus;
wire [temp_w*2-1:0] v2146obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2146 (.l(l[2146*data_w +:data_w]), .r(v2146ibus), .q(v2146obus), .dec(dec[2146]));
wire [data_w*2-1:0] v2147ibus;
wire [temp_w*2-1:0] v2147obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2147 (.l(l[2147*data_w +:data_w]), .r(v2147ibus), .q(v2147obus), .dec(dec[2147]));
wire [data_w*2-1:0] v2148ibus;
wire [temp_w*2-1:0] v2148obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2148 (.l(l[2148*data_w +:data_w]), .r(v2148ibus), .q(v2148obus), .dec(dec[2148]));
wire [data_w*2-1:0] v2149ibus;
wire [temp_w*2-1:0] v2149obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2149 (.l(l[2149*data_w +:data_w]), .r(v2149ibus), .q(v2149obus), .dec(dec[2149]));
wire [data_w*2-1:0] v2150ibus;
wire [temp_w*2-1:0] v2150obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2150 (.l(l[2150*data_w +:data_w]), .r(v2150ibus), .q(v2150obus), .dec(dec[2150]));
wire [data_w*2-1:0] v2151ibus;
wire [temp_w*2-1:0] v2151obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2151 (.l(l[2151*data_w +:data_w]), .r(v2151ibus), .q(v2151obus), .dec(dec[2151]));
wire [data_w*2-1:0] v2152ibus;
wire [temp_w*2-1:0] v2152obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2152 (.l(l[2152*data_w +:data_w]), .r(v2152ibus), .q(v2152obus), .dec(dec[2152]));
wire [data_w*2-1:0] v2153ibus;
wire [temp_w*2-1:0] v2153obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2153 (.l(l[2153*data_w +:data_w]), .r(v2153ibus), .q(v2153obus), .dec(dec[2153]));
wire [data_w*2-1:0] v2154ibus;
wire [temp_w*2-1:0] v2154obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2154 (.l(l[2154*data_w +:data_w]), .r(v2154ibus), .q(v2154obus), .dec(dec[2154]));
wire [data_w*2-1:0] v2155ibus;
wire [temp_w*2-1:0] v2155obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2155 (.l(l[2155*data_w +:data_w]), .r(v2155ibus), .q(v2155obus), .dec(dec[2155]));
wire [data_w*2-1:0] v2156ibus;
wire [temp_w*2-1:0] v2156obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2156 (.l(l[2156*data_w +:data_w]), .r(v2156ibus), .q(v2156obus), .dec(dec[2156]));
wire [data_w*2-1:0] v2157ibus;
wire [temp_w*2-1:0] v2157obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2157 (.l(l[2157*data_w +:data_w]), .r(v2157ibus), .q(v2157obus), .dec(dec[2157]));
wire [data_w*2-1:0] v2158ibus;
wire [temp_w*2-1:0] v2158obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2158 (.l(l[2158*data_w +:data_w]), .r(v2158ibus), .q(v2158obus), .dec(dec[2158]));
wire [data_w*2-1:0] v2159ibus;
wire [temp_w*2-1:0] v2159obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2159 (.l(l[2159*data_w +:data_w]), .r(v2159ibus), .q(v2159obus), .dec(dec[2159]));
wire [data_w*2-1:0] v2160ibus;
wire [temp_w*2-1:0] v2160obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2160 (.l(l[2160*data_w +:data_w]), .r(v2160ibus), .q(v2160obus), .dec(dec[2160]));
wire [data_w*2-1:0] v2161ibus;
wire [temp_w*2-1:0] v2161obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2161 (.l(l[2161*data_w +:data_w]), .r(v2161ibus), .q(v2161obus), .dec(dec[2161]));
wire [data_w*2-1:0] v2162ibus;
wire [temp_w*2-1:0] v2162obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2162 (.l(l[2162*data_w +:data_w]), .r(v2162ibus), .q(v2162obus), .dec(dec[2162]));
wire [data_w*2-1:0] v2163ibus;
wire [temp_w*2-1:0] v2163obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2163 (.l(l[2163*data_w +:data_w]), .r(v2163ibus), .q(v2163obus), .dec(dec[2163]));
wire [data_w*2-1:0] v2164ibus;
wire [temp_w*2-1:0] v2164obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2164 (.l(l[2164*data_w +:data_w]), .r(v2164ibus), .q(v2164obus), .dec(dec[2164]));
wire [data_w*2-1:0] v2165ibus;
wire [temp_w*2-1:0] v2165obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2165 (.l(l[2165*data_w +:data_w]), .r(v2165ibus), .q(v2165obus), .dec(dec[2165]));
wire [data_w*2-1:0] v2166ibus;
wire [temp_w*2-1:0] v2166obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2166 (.l(l[2166*data_w +:data_w]), .r(v2166ibus), .q(v2166obus), .dec(dec[2166]));
wire [data_w*2-1:0] v2167ibus;
wire [temp_w*2-1:0] v2167obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2167 (.l(l[2167*data_w +:data_w]), .r(v2167ibus), .q(v2167obus), .dec(dec[2167]));
wire [data_w*2-1:0] v2168ibus;
wire [temp_w*2-1:0] v2168obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2168 (.l(l[2168*data_w +:data_w]), .r(v2168ibus), .q(v2168obus), .dec(dec[2168]));
wire [data_w*2-1:0] v2169ibus;
wire [temp_w*2-1:0] v2169obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2169 (.l(l[2169*data_w +:data_w]), .r(v2169ibus), .q(v2169obus), .dec(dec[2169]));
wire [data_w*2-1:0] v2170ibus;
wire [temp_w*2-1:0] v2170obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2170 (.l(l[2170*data_w +:data_w]), .r(v2170ibus), .q(v2170obus), .dec(dec[2170]));
wire [data_w*2-1:0] v2171ibus;
wire [temp_w*2-1:0] v2171obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2171 (.l(l[2171*data_w +:data_w]), .r(v2171ibus), .q(v2171obus), .dec(dec[2171]));
wire [data_w*2-1:0] v2172ibus;
wire [temp_w*2-1:0] v2172obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2172 (.l(l[2172*data_w +:data_w]), .r(v2172ibus), .q(v2172obus), .dec(dec[2172]));
wire [data_w*2-1:0] v2173ibus;
wire [temp_w*2-1:0] v2173obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2173 (.l(l[2173*data_w +:data_w]), .r(v2173ibus), .q(v2173obus), .dec(dec[2173]));
wire [data_w*2-1:0] v2174ibus;
wire [temp_w*2-1:0] v2174obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2174 (.l(l[2174*data_w +:data_w]), .r(v2174ibus), .q(v2174obus), .dec(dec[2174]));
wire [data_w*2-1:0] v2175ibus;
wire [temp_w*2-1:0] v2175obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2175 (.l(l[2175*data_w +:data_w]), .r(v2175ibus), .q(v2175obus), .dec(dec[2175]));
wire [data_w*2-1:0] v2176ibus;
wire [temp_w*2-1:0] v2176obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2176 (.l(l[2176*data_w +:data_w]), .r(v2176ibus), .q(v2176obus), .dec(dec[2176]));
wire [data_w*2-1:0] v2177ibus;
wire [temp_w*2-1:0] v2177obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2177 (.l(l[2177*data_w +:data_w]), .r(v2177ibus), .q(v2177obus), .dec(dec[2177]));
wire [data_w*2-1:0] v2178ibus;
wire [temp_w*2-1:0] v2178obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2178 (.l(l[2178*data_w +:data_w]), .r(v2178ibus), .q(v2178obus), .dec(dec[2178]));
wire [data_w*2-1:0] v2179ibus;
wire [temp_w*2-1:0] v2179obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2179 (.l(l[2179*data_w +:data_w]), .r(v2179ibus), .q(v2179obus), .dec(dec[2179]));
wire [data_w*2-1:0] v2180ibus;
wire [temp_w*2-1:0] v2180obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2180 (.l(l[2180*data_w +:data_w]), .r(v2180ibus), .q(v2180obus), .dec(dec[2180]));
wire [data_w*2-1:0] v2181ibus;
wire [temp_w*2-1:0] v2181obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2181 (.l(l[2181*data_w +:data_w]), .r(v2181ibus), .q(v2181obus), .dec(dec[2181]));
wire [data_w*2-1:0] v2182ibus;
wire [temp_w*2-1:0] v2182obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2182 (.l(l[2182*data_w +:data_w]), .r(v2182ibus), .q(v2182obus), .dec(dec[2182]));
wire [data_w*2-1:0] v2183ibus;
wire [temp_w*2-1:0] v2183obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2183 (.l(l[2183*data_w +:data_w]), .r(v2183ibus), .q(v2183obus), .dec(dec[2183]));
wire [data_w*2-1:0] v2184ibus;
wire [temp_w*2-1:0] v2184obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2184 (.l(l[2184*data_w +:data_w]), .r(v2184ibus), .q(v2184obus), .dec(dec[2184]));
wire [data_w*2-1:0] v2185ibus;
wire [temp_w*2-1:0] v2185obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2185 (.l(l[2185*data_w +:data_w]), .r(v2185ibus), .q(v2185obus), .dec(dec[2185]));
wire [data_w*2-1:0] v2186ibus;
wire [temp_w*2-1:0] v2186obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2186 (.l(l[2186*data_w +:data_w]), .r(v2186ibus), .q(v2186obus), .dec(dec[2186]));
wire [data_w*2-1:0] v2187ibus;
wire [temp_w*2-1:0] v2187obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2187 (.l(l[2187*data_w +:data_w]), .r(v2187ibus), .q(v2187obus), .dec(dec[2187]));
wire [data_w*2-1:0] v2188ibus;
wire [temp_w*2-1:0] v2188obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2188 (.l(l[2188*data_w +:data_w]), .r(v2188ibus), .q(v2188obus), .dec(dec[2188]));
wire [data_w*2-1:0] v2189ibus;
wire [temp_w*2-1:0] v2189obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2189 (.l(l[2189*data_w +:data_w]), .r(v2189ibus), .q(v2189obus), .dec(dec[2189]));
wire [data_w*2-1:0] v2190ibus;
wire [temp_w*2-1:0] v2190obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2190 (.l(l[2190*data_w +:data_w]), .r(v2190ibus), .q(v2190obus), .dec(dec[2190]));
wire [data_w*2-1:0] v2191ibus;
wire [temp_w*2-1:0] v2191obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2191 (.l(l[2191*data_w +:data_w]), .r(v2191ibus), .q(v2191obus), .dec(dec[2191]));
wire [data_w*2-1:0] v2192ibus;
wire [temp_w*2-1:0] v2192obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2192 (.l(l[2192*data_w +:data_w]), .r(v2192ibus), .q(v2192obus), .dec(dec[2192]));
wire [data_w*2-1:0] v2193ibus;
wire [temp_w*2-1:0] v2193obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2193 (.l(l[2193*data_w +:data_w]), .r(v2193ibus), .q(v2193obus), .dec(dec[2193]));
wire [data_w*2-1:0] v2194ibus;
wire [temp_w*2-1:0] v2194obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2194 (.l(l[2194*data_w +:data_w]), .r(v2194ibus), .q(v2194obus), .dec(dec[2194]));
wire [data_w*2-1:0] v2195ibus;
wire [temp_w*2-1:0] v2195obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2195 (.l(l[2195*data_w +:data_w]), .r(v2195ibus), .q(v2195obus), .dec(dec[2195]));
wire [data_w*2-1:0] v2196ibus;
wire [temp_w*2-1:0] v2196obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2196 (.l(l[2196*data_w +:data_w]), .r(v2196ibus), .q(v2196obus), .dec(dec[2196]));
wire [data_w*2-1:0] v2197ibus;
wire [temp_w*2-1:0] v2197obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2197 (.l(l[2197*data_w +:data_w]), .r(v2197ibus), .q(v2197obus), .dec(dec[2197]));
wire [data_w*2-1:0] v2198ibus;
wire [temp_w*2-1:0] v2198obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2198 (.l(l[2198*data_w +:data_w]), .r(v2198ibus), .q(v2198obus), .dec(dec[2198]));
wire [data_w*2-1:0] v2199ibus;
wire [temp_w*2-1:0] v2199obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2199 (.l(l[2199*data_w +:data_w]), .r(v2199ibus), .q(v2199obus), .dec(dec[2199]));
wire [data_w*2-1:0] v2200ibus;
wire [temp_w*2-1:0] v2200obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2200 (.l(l[2200*data_w +:data_w]), .r(v2200ibus), .q(v2200obus), .dec(dec[2200]));
wire [data_w*2-1:0] v2201ibus;
wire [temp_w*2-1:0] v2201obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2201 (.l(l[2201*data_w +:data_w]), .r(v2201ibus), .q(v2201obus), .dec(dec[2201]));
wire [data_w*2-1:0] v2202ibus;
wire [temp_w*2-1:0] v2202obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2202 (.l(l[2202*data_w +:data_w]), .r(v2202ibus), .q(v2202obus), .dec(dec[2202]));
wire [data_w*2-1:0] v2203ibus;
wire [temp_w*2-1:0] v2203obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2203 (.l(l[2203*data_w +:data_w]), .r(v2203ibus), .q(v2203obus), .dec(dec[2203]));
wire [data_w*2-1:0] v2204ibus;
wire [temp_w*2-1:0] v2204obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2204 (.l(l[2204*data_w +:data_w]), .r(v2204ibus), .q(v2204obus), .dec(dec[2204]));
wire [data_w*2-1:0] v2205ibus;
wire [temp_w*2-1:0] v2205obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2205 (.l(l[2205*data_w +:data_w]), .r(v2205ibus), .q(v2205obus), .dec(dec[2205]));
wire [data_w*2-1:0] v2206ibus;
wire [temp_w*2-1:0] v2206obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2206 (.l(l[2206*data_w +:data_w]), .r(v2206ibus), .q(v2206obus), .dec(dec[2206]));
wire [data_w*2-1:0] v2207ibus;
wire [temp_w*2-1:0] v2207obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2207 (.l(l[2207*data_w +:data_w]), .r(v2207ibus), .q(v2207obus), .dec(dec[2207]));
wire [data_w*2-1:0] v2208ibus;
wire [temp_w*2-1:0] v2208obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2208 (.l(l[2208*data_w +:data_w]), .r(v2208ibus), .q(v2208obus), .dec(dec[2208]));
wire [data_w*2-1:0] v2209ibus;
wire [temp_w*2-1:0] v2209obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2209 (.l(l[2209*data_w +:data_w]), .r(v2209ibus), .q(v2209obus), .dec(dec[2209]));
wire [data_w*2-1:0] v2210ibus;
wire [temp_w*2-1:0] v2210obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2210 (.l(l[2210*data_w +:data_w]), .r(v2210ibus), .q(v2210obus), .dec(dec[2210]));
wire [data_w*2-1:0] v2211ibus;
wire [temp_w*2-1:0] v2211obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2211 (.l(l[2211*data_w +:data_w]), .r(v2211ibus), .q(v2211obus), .dec(dec[2211]));
wire [data_w*2-1:0] v2212ibus;
wire [temp_w*2-1:0] v2212obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2212 (.l(l[2212*data_w +:data_w]), .r(v2212ibus), .q(v2212obus), .dec(dec[2212]));
wire [data_w*2-1:0] v2213ibus;
wire [temp_w*2-1:0] v2213obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2213 (.l(l[2213*data_w +:data_w]), .r(v2213ibus), .q(v2213obus), .dec(dec[2213]));
wire [data_w*2-1:0] v2214ibus;
wire [temp_w*2-1:0] v2214obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2214 (.l(l[2214*data_w +:data_w]), .r(v2214ibus), .q(v2214obus), .dec(dec[2214]));
wire [data_w*2-1:0] v2215ibus;
wire [temp_w*2-1:0] v2215obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2215 (.l(l[2215*data_w +:data_w]), .r(v2215ibus), .q(v2215obus), .dec(dec[2215]));
wire [data_w*2-1:0] v2216ibus;
wire [temp_w*2-1:0] v2216obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2216 (.l(l[2216*data_w +:data_w]), .r(v2216ibus), .q(v2216obus), .dec(dec[2216]));
wire [data_w*2-1:0] v2217ibus;
wire [temp_w*2-1:0] v2217obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2217 (.l(l[2217*data_w +:data_w]), .r(v2217ibus), .q(v2217obus), .dec(dec[2217]));
wire [data_w*2-1:0] v2218ibus;
wire [temp_w*2-1:0] v2218obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2218 (.l(l[2218*data_w +:data_w]), .r(v2218ibus), .q(v2218obus), .dec(dec[2218]));
wire [data_w*2-1:0] v2219ibus;
wire [temp_w*2-1:0] v2219obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2219 (.l(l[2219*data_w +:data_w]), .r(v2219ibus), .q(v2219obus), .dec(dec[2219]));
wire [data_w*2-1:0] v2220ibus;
wire [temp_w*2-1:0] v2220obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2220 (.l(l[2220*data_w +:data_w]), .r(v2220ibus), .q(v2220obus), .dec(dec[2220]));
wire [data_w*2-1:0] v2221ibus;
wire [temp_w*2-1:0] v2221obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2221 (.l(l[2221*data_w +:data_w]), .r(v2221ibus), .q(v2221obus), .dec(dec[2221]));
wire [data_w*2-1:0] v2222ibus;
wire [temp_w*2-1:0] v2222obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2222 (.l(l[2222*data_w +:data_w]), .r(v2222ibus), .q(v2222obus), .dec(dec[2222]));
wire [data_w*2-1:0] v2223ibus;
wire [temp_w*2-1:0] v2223obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2223 (.l(l[2223*data_w +:data_w]), .r(v2223ibus), .q(v2223obus), .dec(dec[2223]));
wire [data_w*2-1:0] v2224ibus;
wire [temp_w*2-1:0] v2224obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2224 (.l(l[2224*data_w +:data_w]), .r(v2224ibus), .q(v2224obus), .dec(dec[2224]));
wire [data_w*2-1:0] v2225ibus;
wire [temp_w*2-1:0] v2225obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2225 (.l(l[2225*data_w +:data_w]), .r(v2225ibus), .q(v2225obus), .dec(dec[2225]));
wire [data_w*2-1:0] v2226ibus;
wire [temp_w*2-1:0] v2226obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2226 (.l(l[2226*data_w +:data_w]), .r(v2226ibus), .q(v2226obus), .dec(dec[2226]));
wire [data_w*2-1:0] v2227ibus;
wire [temp_w*2-1:0] v2227obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2227 (.l(l[2227*data_w +:data_w]), .r(v2227ibus), .q(v2227obus), .dec(dec[2227]));
wire [data_w*2-1:0] v2228ibus;
wire [temp_w*2-1:0] v2228obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2228 (.l(l[2228*data_w +:data_w]), .r(v2228ibus), .q(v2228obus), .dec(dec[2228]));
wire [data_w*2-1:0] v2229ibus;
wire [temp_w*2-1:0] v2229obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2229 (.l(l[2229*data_w +:data_w]), .r(v2229ibus), .q(v2229obus), .dec(dec[2229]));
wire [data_w*2-1:0] v2230ibus;
wire [temp_w*2-1:0] v2230obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2230 (.l(l[2230*data_w +:data_w]), .r(v2230ibus), .q(v2230obus), .dec(dec[2230]));
wire [data_w*2-1:0] v2231ibus;
wire [temp_w*2-1:0] v2231obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2231 (.l(l[2231*data_w +:data_w]), .r(v2231ibus), .q(v2231obus), .dec(dec[2231]));
wire [data_w*2-1:0] v2232ibus;
wire [temp_w*2-1:0] v2232obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2232 (.l(l[2232*data_w +:data_w]), .r(v2232ibus), .q(v2232obus), .dec(dec[2232]));
wire [data_w*2-1:0] v2233ibus;
wire [temp_w*2-1:0] v2233obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2233 (.l(l[2233*data_w +:data_w]), .r(v2233ibus), .q(v2233obus), .dec(dec[2233]));
wire [data_w*2-1:0] v2234ibus;
wire [temp_w*2-1:0] v2234obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2234 (.l(l[2234*data_w +:data_w]), .r(v2234ibus), .q(v2234obus), .dec(dec[2234]));
wire [data_w*2-1:0] v2235ibus;
wire [temp_w*2-1:0] v2235obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2235 (.l(l[2235*data_w +:data_w]), .r(v2235ibus), .q(v2235obus), .dec(dec[2235]));
wire [data_w*2-1:0] v2236ibus;
wire [temp_w*2-1:0] v2236obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2236 (.l(l[2236*data_w +:data_w]), .r(v2236ibus), .q(v2236obus), .dec(dec[2236]));
wire [data_w*2-1:0] v2237ibus;
wire [temp_w*2-1:0] v2237obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2237 (.l(l[2237*data_w +:data_w]), .r(v2237ibus), .q(v2237obus), .dec(dec[2237]));
wire [data_w*2-1:0] v2238ibus;
wire [temp_w*2-1:0] v2238obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2238 (.l(l[2238*data_w +:data_w]), .r(v2238ibus), .q(v2238obus), .dec(dec[2238]));
wire [data_w*2-1:0] v2239ibus;
wire [temp_w*2-1:0] v2239obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2239 (.l(l[2239*data_w +:data_w]), .r(v2239ibus), .q(v2239obus), .dec(dec[2239]));
wire [data_w*2-1:0] v2240ibus;
wire [temp_w*2-1:0] v2240obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2240 (.l(l[2240*data_w +:data_w]), .r(v2240ibus), .q(v2240obus), .dec(dec[2240]));
wire [data_w*2-1:0] v2241ibus;
wire [temp_w*2-1:0] v2241obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2241 (.l(l[2241*data_w +:data_w]), .r(v2241ibus), .q(v2241obus), .dec(dec[2241]));
wire [data_w*2-1:0] v2242ibus;
wire [temp_w*2-1:0] v2242obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2242 (.l(l[2242*data_w +:data_w]), .r(v2242ibus), .q(v2242obus), .dec(dec[2242]));
wire [data_w*2-1:0] v2243ibus;
wire [temp_w*2-1:0] v2243obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2243 (.l(l[2243*data_w +:data_w]), .r(v2243ibus), .q(v2243obus), .dec(dec[2243]));
wire [data_w*2-1:0] v2244ibus;
wire [temp_w*2-1:0] v2244obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2244 (.l(l[2244*data_w +:data_w]), .r(v2244ibus), .q(v2244obus), .dec(dec[2244]));
wire [data_w*2-1:0] v2245ibus;
wire [temp_w*2-1:0] v2245obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2245 (.l(l[2245*data_w +:data_w]), .r(v2245ibus), .q(v2245obus), .dec(dec[2245]));
wire [data_w*2-1:0] v2246ibus;
wire [temp_w*2-1:0] v2246obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2246 (.l(l[2246*data_w +:data_w]), .r(v2246ibus), .q(v2246obus), .dec(dec[2246]));
wire [data_w*2-1:0] v2247ibus;
wire [temp_w*2-1:0] v2247obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2247 (.l(l[2247*data_w +:data_w]), .r(v2247ibus), .q(v2247obus), .dec(dec[2247]));
wire [data_w*2-1:0] v2248ibus;
wire [temp_w*2-1:0] v2248obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2248 (.l(l[2248*data_w +:data_w]), .r(v2248ibus), .q(v2248obus), .dec(dec[2248]));
wire [data_w*2-1:0] v2249ibus;
wire [temp_w*2-1:0] v2249obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2249 (.l(l[2249*data_w +:data_w]), .r(v2249ibus), .q(v2249obus), .dec(dec[2249]));
wire [data_w*2-1:0] v2250ibus;
wire [temp_w*2-1:0] v2250obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2250 (.l(l[2250*data_w +:data_w]), .r(v2250ibus), .q(v2250obus), .dec(dec[2250]));
wire [data_w*2-1:0] v2251ibus;
wire [temp_w*2-1:0] v2251obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2251 (.l(l[2251*data_w +:data_w]), .r(v2251ibus), .q(v2251obus), .dec(dec[2251]));
wire [data_w*2-1:0] v2252ibus;
wire [temp_w*2-1:0] v2252obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2252 (.l(l[2252*data_w +:data_w]), .r(v2252ibus), .q(v2252obus), .dec(dec[2252]));
wire [data_w*2-1:0] v2253ibus;
wire [temp_w*2-1:0] v2253obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2253 (.l(l[2253*data_w +:data_w]), .r(v2253ibus), .q(v2253obus), .dec(dec[2253]));
wire [data_w*2-1:0] v2254ibus;
wire [temp_w*2-1:0] v2254obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2254 (.l(l[2254*data_w +:data_w]), .r(v2254ibus), .q(v2254obus), .dec(dec[2254]));
wire [data_w*2-1:0] v2255ibus;
wire [temp_w*2-1:0] v2255obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2255 (.l(l[2255*data_w +:data_w]), .r(v2255ibus), .q(v2255obus), .dec(dec[2255]));
wire [data_w*2-1:0] v2256ibus;
wire [temp_w*2-1:0] v2256obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2256 (.l(l[2256*data_w +:data_w]), .r(v2256ibus), .q(v2256obus), .dec(dec[2256]));
wire [data_w*2-1:0] v2257ibus;
wire [temp_w*2-1:0] v2257obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2257 (.l(l[2257*data_w +:data_w]), .r(v2257ibus), .q(v2257obus), .dec(dec[2257]));
wire [data_w*2-1:0] v2258ibus;
wire [temp_w*2-1:0] v2258obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2258 (.l(l[2258*data_w +:data_w]), .r(v2258ibus), .q(v2258obus), .dec(dec[2258]));
wire [data_w*2-1:0] v2259ibus;
wire [temp_w*2-1:0] v2259obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2259 (.l(l[2259*data_w +:data_w]), .r(v2259ibus), .q(v2259obus), .dec(dec[2259]));
wire [data_w*2-1:0] v2260ibus;
wire [temp_w*2-1:0] v2260obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2260 (.l(l[2260*data_w +:data_w]), .r(v2260ibus), .q(v2260obus), .dec(dec[2260]));
wire [data_w*2-1:0] v2261ibus;
wire [temp_w*2-1:0] v2261obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2261 (.l(l[2261*data_w +:data_w]), .r(v2261ibus), .q(v2261obus), .dec(dec[2261]));
wire [data_w*2-1:0] v2262ibus;
wire [temp_w*2-1:0] v2262obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2262 (.l(l[2262*data_w +:data_w]), .r(v2262ibus), .q(v2262obus), .dec(dec[2262]));
wire [data_w*2-1:0] v2263ibus;
wire [temp_w*2-1:0] v2263obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2263 (.l(l[2263*data_w +:data_w]), .r(v2263ibus), .q(v2263obus), .dec(dec[2263]));
wire [data_w*2-1:0] v2264ibus;
wire [temp_w*2-1:0] v2264obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2264 (.l(l[2264*data_w +:data_w]), .r(v2264ibus), .q(v2264obus), .dec(dec[2264]));
wire [data_w*2-1:0] v2265ibus;
wire [temp_w*2-1:0] v2265obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2265 (.l(l[2265*data_w +:data_w]), .r(v2265ibus), .q(v2265obus), .dec(dec[2265]));
wire [data_w*2-1:0] v2266ibus;
wire [temp_w*2-1:0] v2266obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2266 (.l(l[2266*data_w +:data_w]), .r(v2266ibus), .q(v2266obus), .dec(dec[2266]));
wire [data_w*2-1:0] v2267ibus;
wire [temp_w*2-1:0] v2267obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2267 (.l(l[2267*data_w +:data_w]), .r(v2267ibus), .q(v2267obus), .dec(dec[2267]));
wire [data_w*2-1:0] v2268ibus;
wire [temp_w*2-1:0] v2268obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2268 (.l(l[2268*data_w +:data_w]), .r(v2268ibus), .q(v2268obus), .dec(dec[2268]));
wire [data_w*2-1:0] v2269ibus;
wire [temp_w*2-1:0] v2269obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2269 (.l(l[2269*data_w +:data_w]), .r(v2269ibus), .q(v2269obus), .dec(dec[2269]));
wire [data_w*2-1:0] v2270ibus;
wire [temp_w*2-1:0] v2270obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2270 (.l(l[2270*data_w +:data_w]), .r(v2270ibus), .q(v2270obus), .dec(dec[2270]));
wire [data_w*2-1:0] v2271ibus;
wire [temp_w*2-1:0] v2271obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2271 (.l(l[2271*data_w +:data_w]), .r(v2271ibus), .q(v2271obus), .dec(dec[2271]));
wire [data_w*2-1:0] v2272ibus;
wire [temp_w*2-1:0] v2272obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2272 (.l(l[2272*data_w +:data_w]), .r(v2272ibus), .q(v2272obus), .dec(dec[2272]));
wire [data_w*2-1:0] v2273ibus;
wire [temp_w*2-1:0] v2273obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2273 (.l(l[2273*data_w +:data_w]), .r(v2273ibus), .q(v2273obus), .dec(dec[2273]));
wire [data_w*2-1:0] v2274ibus;
wire [temp_w*2-1:0] v2274obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2274 (.l(l[2274*data_w +:data_w]), .r(v2274ibus), .q(v2274obus), .dec(dec[2274]));
wire [data_w*2-1:0] v2275ibus;
wire [temp_w*2-1:0] v2275obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2275 (.l(l[2275*data_w +:data_w]), .r(v2275ibus), .q(v2275obus), .dec(dec[2275]));
wire [data_w*2-1:0] v2276ibus;
wire [temp_w*2-1:0] v2276obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2276 (.l(l[2276*data_w +:data_w]), .r(v2276ibus), .q(v2276obus), .dec(dec[2276]));
wire [data_w*2-1:0] v2277ibus;
wire [temp_w*2-1:0] v2277obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2277 (.l(l[2277*data_w +:data_w]), .r(v2277ibus), .q(v2277obus), .dec(dec[2277]));
wire [data_w*2-1:0] v2278ibus;
wire [temp_w*2-1:0] v2278obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2278 (.l(l[2278*data_w +:data_w]), .r(v2278ibus), .q(v2278obus), .dec(dec[2278]));
wire [data_w*2-1:0] v2279ibus;
wire [temp_w*2-1:0] v2279obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2279 (.l(l[2279*data_w +:data_w]), .r(v2279ibus), .q(v2279obus), .dec(dec[2279]));
wire [data_w*2-1:0] v2280ibus;
wire [temp_w*2-1:0] v2280obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2280 (.l(l[2280*data_w +:data_w]), .r(v2280ibus), .q(v2280obus), .dec(dec[2280]));
wire [data_w*2-1:0] v2281ibus;
wire [temp_w*2-1:0] v2281obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2281 (.l(l[2281*data_w +:data_w]), .r(v2281ibus), .q(v2281obus), .dec(dec[2281]));
wire [data_w*2-1:0] v2282ibus;
wire [temp_w*2-1:0] v2282obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2282 (.l(l[2282*data_w +:data_w]), .r(v2282ibus), .q(v2282obus), .dec(dec[2282]));
wire [data_w*2-1:0] v2283ibus;
wire [temp_w*2-1:0] v2283obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2283 (.l(l[2283*data_w +:data_w]), .r(v2283ibus), .q(v2283obus), .dec(dec[2283]));
wire [data_w*2-1:0] v2284ibus;
wire [temp_w*2-1:0] v2284obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2284 (.l(l[2284*data_w +:data_w]), .r(v2284ibus), .q(v2284obus), .dec(dec[2284]));
wire [data_w*2-1:0] v2285ibus;
wire [temp_w*2-1:0] v2285obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2285 (.l(l[2285*data_w +:data_w]), .r(v2285ibus), .q(v2285obus), .dec(dec[2285]));
wire [data_w*2-1:0] v2286ibus;
wire [temp_w*2-1:0] v2286obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2286 (.l(l[2286*data_w +:data_w]), .r(v2286ibus), .q(v2286obus), .dec(dec[2286]));
wire [data_w*2-1:0] v2287ibus;
wire [temp_w*2-1:0] v2287obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2287 (.l(l[2287*data_w +:data_w]), .r(v2287ibus), .q(v2287obus), .dec(dec[2287]));
wire [data_w*2-1:0] v2288ibus;
wire [temp_w*2-1:0] v2288obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2288 (.l(l[2288*data_w +:data_w]), .r(v2288ibus), .q(v2288obus), .dec(dec[2288]));
wire [data_w*2-1:0] v2289ibus;
wire [temp_w*2-1:0] v2289obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2289 (.l(l[2289*data_w +:data_w]), .r(v2289ibus), .q(v2289obus), .dec(dec[2289]));
wire [data_w*2-1:0] v2290ibus;
wire [temp_w*2-1:0] v2290obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2290 (.l(l[2290*data_w +:data_w]), .r(v2290ibus), .q(v2290obus), .dec(dec[2290]));
wire [data_w*2-1:0] v2291ibus;
wire [temp_w*2-1:0] v2291obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2291 (.l(l[2291*data_w +:data_w]), .r(v2291ibus), .q(v2291obus), .dec(dec[2291]));
wire [data_w*2-1:0] v2292ibus;
wire [temp_w*2-1:0] v2292obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2292 (.l(l[2292*data_w +:data_w]), .r(v2292ibus), .q(v2292obus), .dec(dec[2292]));
wire [data_w*2-1:0] v2293ibus;
wire [temp_w*2-1:0] v2293obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2293 (.l(l[2293*data_w +:data_w]), .r(v2293ibus), .q(v2293obus), .dec(dec[2293]));
wire [data_w*2-1:0] v2294ibus;
wire [temp_w*2-1:0] v2294obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2294 (.l(l[2294*data_w +:data_w]), .r(v2294ibus), .q(v2294obus), .dec(dec[2294]));
wire [data_w*2-1:0] v2295ibus;
wire [temp_w*2-1:0] v2295obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2295 (.l(l[2295*data_w +:data_w]), .r(v2295ibus), .q(v2295obus), .dec(dec[2295]));
wire [data_w*2-1:0] v2296ibus;
wire [temp_w*2-1:0] v2296obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2296 (.l(l[2296*data_w +:data_w]), .r(v2296ibus), .q(v2296obus), .dec(dec[2296]));
wire [data_w*2-1:0] v2297ibus;
wire [temp_w*2-1:0] v2297obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2297 (.l(l[2297*data_w +:data_w]), .r(v2297ibus), .q(v2297obus), .dec(dec[2297]));
wire [data_w*2-1:0] v2298ibus;
wire [temp_w*2-1:0] v2298obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2298 (.l(l[2298*data_w +:data_w]), .r(v2298ibus), .q(v2298obus), .dec(dec[2298]));
wire [data_w*2-1:0] v2299ibus;
wire [temp_w*2-1:0] v2299obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2299 (.l(l[2299*data_w +:data_w]), .r(v2299ibus), .q(v2299obus), .dec(dec[2299]));
wire [data_w*2-1:0] v2300ibus;
wire [temp_w*2-1:0] v2300obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2300 (.l(l[2300*data_w +:data_w]), .r(v2300ibus), .q(v2300obus), .dec(dec[2300]));
wire [data_w*2-1:0] v2301ibus;
wire [temp_w*2-1:0] v2301obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2301 (.l(l[2301*data_w +:data_w]), .r(v2301ibus), .q(v2301obus), .dec(dec[2301]));
wire [data_w*2-1:0] v2302ibus;
wire [temp_w*2-1:0] v2302obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2302 (.l(l[2302*data_w +:data_w]), .r(v2302ibus), .q(v2302obus), .dec(dec[2302]));
wire [data_w*2-1:0] v2303ibus;
wire [temp_w*2-1:0] v2303obus;
vnu #(.data_w(data_w), .D(2), .ext_w(ext_w)) VNU2303 (.l(l[2303*data_w +:data_w]), .r(v2303ibus), .q(v2303obus), .dec(dec[2303]));
assign c0ibus[temp_w*0 +:temp_w] = v190obus[temp_w*0 +:temp_w];
assign v190ibus[data_w*0 +:data_w] = c0obus[data_w*0 +:data_w];
assign c0ibus[temp_w*1 +:temp_w] = v265obus[temp_w*0 +:temp_w];
assign v265ibus[data_w*0 +:data_w] = c0obus[data_w*1 +:data_w];
assign c0ibus[temp_w*2 +:temp_w] = v823obus[temp_w*0 +:temp_w];
assign v823ibus[data_w*0 +:data_w] = c0obus[data_w*2 +:data_w];
assign c0ibus[temp_w*3 +:temp_w] = v947obus[temp_w*0 +:temp_w];
assign v947ibus[data_w*0 +:data_w] = c0obus[data_w*3 +:data_w];
assign c0ibus[temp_w*4 +:temp_w] = v1159obus[temp_w*0 +:temp_w];
assign v1159ibus[data_w*0 +:data_w] = c0obus[data_w*4 +:data_w];
assign c0ibus[temp_w*5 +:temp_w] = v1248obus[temp_w*0 +:temp_w];
assign v1248ibus[data_w*0 +:data_w] = c0obus[data_w*5 +:data_w];
assign c1ibus[temp_w*0 +:temp_w] = v191obus[temp_w*0 +:temp_w];
assign v191ibus[data_w*0 +:data_w] = c1obus[data_w*0 +:data_w];
assign c1ibus[temp_w*1 +:temp_w] = v266obus[temp_w*0 +:temp_w];
assign v266ibus[data_w*0 +:data_w] = c1obus[data_w*1 +:data_w];
assign c1ibus[temp_w*2 +:temp_w] = v824obus[temp_w*0 +:temp_w];
assign v824ibus[data_w*0 +:data_w] = c1obus[data_w*2 +:data_w];
assign c1ibus[temp_w*3 +:temp_w] = v948obus[temp_w*0 +:temp_w];
assign v948ibus[data_w*0 +:data_w] = c1obus[data_w*3 +:data_w];
assign c1ibus[temp_w*4 +:temp_w] = v1160obus[temp_w*0 +:temp_w];
assign v1160ibus[data_w*0 +:data_w] = c1obus[data_w*4 +:data_w];
assign c1ibus[temp_w*5 +:temp_w] = v1249obus[temp_w*0 +:temp_w];
assign v1249ibus[data_w*0 +:data_w] = c1obus[data_w*5 +:data_w];
assign c2ibus[temp_w*0 +:temp_w] = v96obus[temp_w*0 +:temp_w];
assign v96ibus[data_w*0 +:data_w] = c2obus[data_w*0 +:data_w];
assign c2ibus[temp_w*1 +:temp_w] = v267obus[temp_w*0 +:temp_w];
assign v267ibus[data_w*0 +:data_w] = c2obus[data_w*1 +:data_w];
assign c2ibus[temp_w*2 +:temp_w] = v825obus[temp_w*0 +:temp_w];
assign v825ibus[data_w*0 +:data_w] = c2obus[data_w*2 +:data_w];
assign c2ibus[temp_w*3 +:temp_w] = v949obus[temp_w*0 +:temp_w];
assign v949ibus[data_w*0 +:data_w] = c2obus[data_w*3 +:data_w];
assign c2ibus[temp_w*4 +:temp_w] = v1161obus[temp_w*0 +:temp_w];
assign v1161ibus[data_w*0 +:data_w] = c2obus[data_w*4 +:data_w];
assign c2ibus[temp_w*5 +:temp_w] = v1250obus[temp_w*0 +:temp_w];
assign v1250ibus[data_w*0 +:data_w] = c2obus[data_w*5 +:data_w];
assign c3ibus[temp_w*0 +:temp_w] = v97obus[temp_w*0 +:temp_w];
assign v97ibus[data_w*0 +:data_w] = c3obus[data_w*0 +:data_w];
assign c3ibus[temp_w*1 +:temp_w] = v268obus[temp_w*0 +:temp_w];
assign v268ibus[data_w*0 +:data_w] = c3obus[data_w*1 +:data_w];
assign c3ibus[temp_w*2 +:temp_w] = v826obus[temp_w*0 +:temp_w];
assign v826ibus[data_w*0 +:data_w] = c3obus[data_w*2 +:data_w];
assign c3ibus[temp_w*3 +:temp_w] = v950obus[temp_w*0 +:temp_w];
assign v950ibus[data_w*0 +:data_w] = c3obus[data_w*3 +:data_w];
assign c3ibus[temp_w*4 +:temp_w] = v1162obus[temp_w*0 +:temp_w];
assign v1162ibus[data_w*0 +:data_w] = c3obus[data_w*4 +:data_w];
assign c3ibus[temp_w*5 +:temp_w] = v1251obus[temp_w*0 +:temp_w];
assign v1251ibus[data_w*0 +:data_w] = c3obus[data_w*5 +:data_w];
assign c4ibus[temp_w*0 +:temp_w] = v98obus[temp_w*0 +:temp_w];
assign v98ibus[data_w*0 +:data_w] = c4obus[data_w*0 +:data_w];
assign c4ibus[temp_w*1 +:temp_w] = v269obus[temp_w*0 +:temp_w];
assign v269ibus[data_w*0 +:data_w] = c4obus[data_w*1 +:data_w];
assign c4ibus[temp_w*2 +:temp_w] = v827obus[temp_w*0 +:temp_w];
assign v827ibus[data_w*0 +:data_w] = c4obus[data_w*2 +:data_w];
assign c4ibus[temp_w*3 +:temp_w] = v951obus[temp_w*0 +:temp_w];
assign v951ibus[data_w*0 +:data_w] = c4obus[data_w*3 +:data_w];
assign c4ibus[temp_w*4 +:temp_w] = v1163obus[temp_w*0 +:temp_w];
assign v1163ibus[data_w*0 +:data_w] = c4obus[data_w*4 +:data_w];
assign c4ibus[temp_w*5 +:temp_w] = v1252obus[temp_w*0 +:temp_w];
assign v1252ibus[data_w*0 +:data_w] = c4obus[data_w*5 +:data_w];
assign c5ibus[temp_w*0 +:temp_w] = v99obus[temp_w*0 +:temp_w];
assign v99ibus[data_w*0 +:data_w] = c5obus[data_w*0 +:data_w];
assign c5ibus[temp_w*1 +:temp_w] = v270obus[temp_w*0 +:temp_w];
assign v270ibus[data_w*0 +:data_w] = c5obus[data_w*1 +:data_w];
assign c5ibus[temp_w*2 +:temp_w] = v828obus[temp_w*0 +:temp_w];
assign v828ibus[data_w*0 +:data_w] = c5obus[data_w*2 +:data_w];
assign c5ibus[temp_w*3 +:temp_w] = v952obus[temp_w*0 +:temp_w];
assign v952ibus[data_w*0 +:data_w] = c5obus[data_w*3 +:data_w];
assign c5ibus[temp_w*4 +:temp_w] = v1164obus[temp_w*0 +:temp_w];
assign v1164ibus[data_w*0 +:data_w] = c5obus[data_w*4 +:data_w];
assign c5ibus[temp_w*5 +:temp_w] = v1253obus[temp_w*0 +:temp_w];
assign v1253ibus[data_w*0 +:data_w] = c5obus[data_w*5 +:data_w];
assign c6ibus[temp_w*0 +:temp_w] = v100obus[temp_w*0 +:temp_w];
assign v100ibus[data_w*0 +:data_w] = c6obus[data_w*0 +:data_w];
assign c6ibus[temp_w*1 +:temp_w] = v271obus[temp_w*0 +:temp_w];
assign v271ibus[data_w*0 +:data_w] = c6obus[data_w*1 +:data_w];
assign c6ibus[temp_w*2 +:temp_w] = v829obus[temp_w*0 +:temp_w];
assign v829ibus[data_w*0 +:data_w] = c6obus[data_w*2 +:data_w];
assign c6ibus[temp_w*3 +:temp_w] = v953obus[temp_w*0 +:temp_w];
assign v953ibus[data_w*0 +:data_w] = c6obus[data_w*3 +:data_w];
assign c6ibus[temp_w*4 +:temp_w] = v1165obus[temp_w*0 +:temp_w];
assign v1165ibus[data_w*0 +:data_w] = c6obus[data_w*4 +:data_w];
assign c6ibus[temp_w*5 +:temp_w] = v1254obus[temp_w*0 +:temp_w];
assign v1254ibus[data_w*0 +:data_w] = c6obus[data_w*5 +:data_w];
assign c7ibus[temp_w*0 +:temp_w] = v101obus[temp_w*0 +:temp_w];
assign v101ibus[data_w*0 +:data_w] = c7obus[data_w*0 +:data_w];
assign c7ibus[temp_w*1 +:temp_w] = v272obus[temp_w*0 +:temp_w];
assign v272ibus[data_w*0 +:data_w] = c7obus[data_w*1 +:data_w];
assign c7ibus[temp_w*2 +:temp_w] = v830obus[temp_w*0 +:temp_w];
assign v830ibus[data_w*0 +:data_w] = c7obus[data_w*2 +:data_w];
assign c7ibus[temp_w*3 +:temp_w] = v954obus[temp_w*0 +:temp_w];
assign v954ibus[data_w*0 +:data_w] = c7obus[data_w*3 +:data_w];
assign c7ibus[temp_w*4 +:temp_w] = v1166obus[temp_w*0 +:temp_w];
assign v1166ibus[data_w*0 +:data_w] = c7obus[data_w*4 +:data_w];
assign c7ibus[temp_w*5 +:temp_w] = v1255obus[temp_w*0 +:temp_w];
assign v1255ibus[data_w*0 +:data_w] = c7obus[data_w*5 +:data_w];
assign c8ibus[temp_w*0 +:temp_w] = v102obus[temp_w*0 +:temp_w];
assign v102ibus[data_w*0 +:data_w] = c8obus[data_w*0 +:data_w];
assign c8ibus[temp_w*1 +:temp_w] = v273obus[temp_w*0 +:temp_w];
assign v273ibus[data_w*0 +:data_w] = c8obus[data_w*1 +:data_w];
assign c8ibus[temp_w*2 +:temp_w] = v831obus[temp_w*0 +:temp_w];
assign v831ibus[data_w*0 +:data_w] = c8obus[data_w*2 +:data_w];
assign c8ibus[temp_w*3 +:temp_w] = v955obus[temp_w*0 +:temp_w];
assign v955ibus[data_w*0 +:data_w] = c8obus[data_w*3 +:data_w];
assign c8ibus[temp_w*4 +:temp_w] = v1167obus[temp_w*0 +:temp_w];
assign v1167ibus[data_w*0 +:data_w] = c8obus[data_w*4 +:data_w];
assign c8ibus[temp_w*5 +:temp_w] = v1256obus[temp_w*0 +:temp_w];
assign v1256ibus[data_w*0 +:data_w] = c8obus[data_w*5 +:data_w];
assign c9ibus[temp_w*0 +:temp_w] = v103obus[temp_w*0 +:temp_w];
assign v103ibus[data_w*0 +:data_w] = c9obus[data_w*0 +:data_w];
assign c9ibus[temp_w*1 +:temp_w] = v274obus[temp_w*0 +:temp_w];
assign v274ibus[data_w*0 +:data_w] = c9obus[data_w*1 +:data_w];
assign c9ibus[temp_w*2 +:temp_w] = v832obus[temp_w*0 +:temp_w];
assign v832ibus[data_w*0 +:data_w] = c9obus[data_w*2 +:data_w];
assign c9ibus[temp_w*3 +:temp_w] = v956obus[temp_w*0 +:temp_w];
assign v956ibus[data_w*0 +:data_w] = c9obus[data_w*3 +:data_w];
assign c9ibus[temp_w*4 +:temp_w] = v1168obus[temp_w*0 +:temp_w];
assign v1168ibus[data_w*0 +:data_w] = c9obus[data_w*4 +:data_w];
assign c9ibus[temp_w*5 +:temp_w] = v1257obus[temp_w*0 +:temp_w];
assign v1257ibus[data_w*0 +:data_w] = c9obus[data_w*5 +:data_w];
assign c10ibus[temp_w*0 +:temp_w] = v104obus[temp_w*0 +:temp_w];
assign v104ibus[data_w*0 +:data_w] = c10obus[data_w*0 +:data_w];
assign c10ibus[temp_w*1 +:temp_w] = v275obus[temp_w*0 +:temp_w];
assign v275ibus[data_w*0 +:data_w] = c10obus[data_w*1 +:data_w];
assign c10ibus[temp_w*2 +:temp_w] = v833obus[temp_w*0 +:temp_w];
assign v833ibus[data_w*0 +:data_w] = c10obus[data_w*2 +:data_w];
assign c10ibus[temp_w*3 +:temp_w] = v957obus[temp_w*0 +:temp_w];
assign v957ibus[data_w*0 +:data_w] = c10obus[data_w*3 +:data_w];
assign c10ibus[temp_w*4 +:temp_w] = v1169obus[temp_w*0 +:temp_w];
assign v1169ibus[data_w*0 +:data_w] = c10obus[data_w*4 +:data_w];
assign c10ibus[temp_w*5 +:temp_w] = v1258obus[temp_w*0 +:temp_w];
assign v1258ibus[data_w*0 +:data_w] = c10obus[data_w*5 +:data_w];
assign c11ibus[temp_w*0 +:temp_w] = v105obus[temp_w*0 +:temp_w];
assign v105ibus[data_w*0 +:data_w] = c11obus[data_w*0 +:data_w];
assign c11ibus[temp_w*1 +:temp_w] = v276obus[temp_w*0 +:temp_w];
assign v276ibus[data_w*0 +:data_w] = c11obus[data_w*1 +:data_w];
assign c11ibus[temp_w*2 +:temp_w] = v834obus[temp_w*0 +:temp_w];
assign v834ibus[data_w*0 +:data_w] = c11obus[data_w*2 +:data_w];
assign c11ibus[temp_w*3 +:temp_w] = v958obus[temp_w*0 +:temp_w];
assign v958ibus[data_w*0 +:data_w] = c11obus[data_w*3 +:data_w];
assign c11ibus[temp_w*4 +:temp_w] = v1170obus[temp_w*0 +:temp_w];
assign v1170ibus[data_w*0 +:data_w] = c11obus[data_w*4 +:data_w];
assign c11ibus[temp_w*5 +:temp_w] = v1259obus[temp_w*0 +:temp_w];
assign v1259ibus[data_w*0 +:data_w] = c11obus[data_w*5 +:data_w];
assign c12ibus[temp_w*0 +:temp_w] = v106obus[temp_w*0 +:temp_w];
assign v106ibus[data_w*0 +:data_w] = c12obus[data_w*0 +:data_w];
assign c12ibus[temp_w*1 +:temp_w] = v277obus[temp_w*0 +:temp_w];
assign v277ibus[data_w*0 +:data_w] = c12obus[data_w*1 +:data_w];
assign c12ibus[temp_w*2 +:temp_w] = v835obus[temp_w*0 +:temp_w];
assign v835ibus[data_w*0 +:data_w] = c12obus[data_w*2 +:data_w];
assign c12ibus[temp_w*3 +:temp_w] = v959obus[temp_w*0 +:temp_w];
assign v959ibus[data_w*0 +:data_w] = c12obus[data_w*3 +:data_w];
assign c12ibus[temp_w*4 +:temp_w] = v1171obus[temp_w*0 +:temp_w];
assign v1171ibus[data_w*0 +:data_w] = c12obus[data_w*4 +:data_w];
assign c12ibus[temp_w*5 +:temp_w] = v1260obus[temp_w*0 +:temp_w];
assign v1260ibus[data_w*0 +:data_w] = c12obus[data_w*5 +:data_w];
assign c13ibus[temp_w*0 +:temp_w] = v107obus[temp_w*0 +:temp_w];
assign v107ibus[data_w*0 +:data_w] = c13obus[data_w*0 +:data_w];
assign c13ibus[temp_w*1 +:temp_w] = v278obus[temp_w*0 +:temp_w];
assign v278ibus[data_w*0 +:data_w] = c13obus[data_w*1 +:data_w];
assign c13ibus[temp_w*2 +:temp_w] = v836obus[temp_w*0 +:temp_w];
assign v836ibus[data_w*0 +:data_w] = c13obus[data_w*2 +:data_w];
assign c13ibus[temp_w*3 +:temp_w] = v864obus[temp_w*0 +:temp_w];
assign v864ibus[data_w*0 +:data_w] = c13obus[data_w*3 +:data_w];
assign c13ibus[temp_w*4 +:temp_w] = v1172obus[temp_w*0 +:temp_w];
assign v1172ibus[data_w*0 +:data_w] = c13obus[data_w*4 +:data_w];
assign c13ibus[temp_w*5 +:temp_w] = v1261obus[temp_w*0 +:temp_w];
assign v1261ibus[data_w*0 +:data_w] = c13obus[data_w*5 +:data_w];
assign c14ibus[temp_w*0 +:temp_w] = v108obus[temp_w*0 +:temp_w];
assign v108ibus[data_w*0 +:data_w] = c14obus[data_w*0 +:data_w];
assign c14ibus[temp_w*1 +:temp_w] = v279obus[temp_w*0 +:temp_w];
assign v279ibus[data_w*0 +:data_w] = c14obus[data_w*1 +:data_w];
assign c14ibus[temp_w*2 +:temp_w] = v837obus[temp_w*0 +:temp_w];
assign v837ibus[data_w*0 +:data_w] = c14obus[data_w*2 +:data_w];
assign c14ibus[temp_w*3 +:temp_w] = v865obus[temp_w*0 +:temp_w];
assign v865ibus[data_w*0 +:data_w] = c14obus[data_w*3 +:data_w];
assign c14ibus[temp_w*4 +:temp_w] = v1173obus[temp_w*0 +:temp_w];
assign v1173ibus[data_w*0 +:data_w] = c14obus[data_w*4 +:data_w];
assign c14ibus[temp_w*5 +:temp_w] = v1262obus[temp_w*0 +:temp_w];
assign v1262ibus[data_w*0 +:data_w] = c14obus[data_w*5 +:data_w];
assign c15ibus[temp_w*0 +:temp_w] = v109obus[temp_w*0 +:temp_w];
assign v109ibus[data_w*0 +:data_w] = c15obus[data_w*0 +:data_w];
assign c15ibus[temp_w*1 +:temp_w] = v280obus[temp_w*0 +:temp_w];
assign v280ibus[data_w*0 +:data_w] = c15obus[data_w*1 +:data_w];
assign c15ibus[temp_w*2 +:temp_w] = v838obus[temp_w*0 +:temp_w];
assign v838ibus[data_w*0 +:data_w] = c15obus[data_w*2 +:data_w];
assign c15ibus[temp_w*3 +:temp_w] = v866obus[temp_w*0 +:temp_w];
assign v866ibus[data_w*0 +:data_w] = c15obus[data_w*3 +:data_w];
assign c15ibus[temp_w*4 +:temp_w] = v1174obus[temp_w*0 +:temp_w];
assign v1174ibus[data_w*0 +:data_w] = c15obus[data_w*4 +:data_w];
assign c15ibus[temp_w*5 +:temp_w] = v1263obus[temp_w*0 +:temp_w];
assign v1263ibus[data_w*0 +:data_w] = c15obus[data_w*5 +:data_w];
assign c16ibus[temp_w*0 +:temp_w] = v110obus[temp_w*0 +:temp_w];
assign v110ibus[data_w*0 +:data_w] = c16obus[data_w*0 +:data_w];
assign c16ibus[temp_w*1 +:temp_w] = v281obus[temp_w*0 +:temp_w];
assign v281ibus[data_w*0 +:data_w] = c16obus[data_w*1 +:data_w];
assign c16ibus[temp_w*2 +:temp_w] = v839obus[temp_w*0 +:temp_w];
assign v839ibus[data_w*0 +:data_w] = c16obus[data_w*2 +:data_w];
assign c16ibus[temp_w*3 +:temp_w] = v867obus[temp_w*0 +:temp_w];
assign v867ibus[data_w*0 +:data_w] = c16obus[data_w*3 +:data_w];
assign c16ibus[temp_w*4 +:temp_w] = v1175obus[temp_w*0 +:temp_w];
assign v1175ibus[data_w*0 +:data_w] = c16obus[data_w*4 +:data_w];
assign c16ibus[temp_w*5 +:temp_w] = v1264obus[temp_w*0 +:temp_w];
assign v1264ibus[data_w*0 +:data_w] = c16obus[data_w*5 +:data_w];
assign c17ibus[temp_w*0 +:temp_w] = v111obus[temp_w*0 +:temp_w];
assign v111ibus[data_w*0 +:data_w] = c17obus[data_w*0 +:data_w];
assign c17ibus[temp_w*1 +:temp_w] = v282obus[temp_w*0 +:temp_w];
assign v282ibus[data_w*0 +:data_w] = c17obus[data_w*1 +:data_w];
assign c17ibus[temp_w*2 +:temp_w] = v840obus[temp_w*0 +:temp_w];
assign v840ibus[data_w*0 +:data_w] = c17obus[data_w*2 +:data_w];
assign c17ibus[temp_w*3 +:temp_w] = v868obus[temp_w*0 +:temp_w];
assign v868ibus[data_w*0 +:data_w] = c17obus[data_w*3 +:data_w];
assign c17ibus[temp_w*4 +:temp_w] = v1176obus[temp_w*0 +:temp_w];
assign v1176ibus[data_w*0 +:data_w] = c17obus[data_w*4 +:data_w];
assign c17ibus[temp_w*5 +:temp_w] = v1265obus[temp_w*0 +:temp_w];
assign v1265ibus[data_w*0 +:data_w] = c17obus[data_w*5 +:data_w];
assign c18ibus[temp_w*0 +:temp_w] = v112obus[temp_w*0 +:temp_w];
assign v112ibus[data_w*0 +:data_w] = c18obus[data_w*0 +:data_w];
assign c18ibus[temp_w*1 +:temp_w] = v283obus[temp_w*0 +:temp_w];
assign v283ibus[data_w*0 +:data_w] = c18obus[data_w*1 +:data_w];
assign c18ibus[temp_w*2 +:temp_w] = v841obus[temp_w*0 +:temp_w];
assign v841ibus[data_w*0 +:data_w] = c18obus[data_w*2 +:data_w];
assign c18ibus[temp_w*3 +:temp_w] = v869obus[temp_w*0 +:temp_w];
assign v869ibus[data_w*0 +:data_w] = c18obus[data_w*3 +:data_w];
assign c18ibus[temp_w*4 +:temp_w] = v1177obus[temp_w*0 +:temp_w];
assign v1177ibus[data_w*0 +:data_w] = c18obus[data_w*4 +:data_w];
assign c18ibus[temp_w*5 +:temp_w] = v1266obus[temp_w*0 +:temp_w];
assign v1266ibus[data_w*0 +:data_w] = c18obus[data_w*5 +:data_w];
assign c19ibus[temp_w*0 +:temp_w] = v113obus[temp_w*0 +:temp_w];
assign v113ibus[data_w*0 +:data_w] = c19obus[data_w*0 +:data_w];
assign c19ibus[temp_w*1 +:temp_w] = v284obus[temp_w*0 +:temp_w];
assign v284ibus[data_w*0 +:data_w] = c19obus[data_w*1 +:data_w];
assign c19ibus[temp_w*2 +:temp_w] = v842obus[temp_w*0 +:temp_w];
assign v842ibus[data_w*0 +:data_w] = c19obus[data_w*2 +:data_w];
assign c19ibus[temp_w*3 +:temp_w] = v870obus[temp_w*0 +:temp_w];
assign v870ibus[data_w*0 +:data_w] = c19obus[data_w*3 +:data_w];
assign c19ibus[temp_w*4 +:temp_w] = v1178obus[temp_w*0 +:temp_w];
assign v1178ibus[data_w*0 +:data_w] = c19obus[data_w*4 +:data_w];
assign c19ibus[temp_w*5 +:temp_w] = v1267obus[temp_w*0 +:temp_w];
assign v1267ibus[data_w*0 +:data_w] = c19obus[data_w*5 +:data_w];
assign c20ibus[temp_w*0 +:temp_w] = v114obus[temp_w*0 +:temp_w];
assign v114ibus[data_w*0 +:data_w] = c20obus[data_w*0 +:data_w];
assign c20ibus[temp_w*1 +:temp_w] = v285obus[temp_w*0 +:temp_w];
assign v285ibus[data_w*0 +:data_w] = c20obus[data_w*1 +:data_w];
assign c20ibus[temp_w*2 +:temp_w] = v843obus[temp_w*0 +:temp_w];
assign v843ibus[data_w*0 +:data_w] = c20obus[data_w*2 +:data_w];
assign c20ibus[temp_w*3 +:temp_w] = v871obus[temp_w*0 +:temp_w];
assign v871ibus[data_w*0 +:data_w] = c20obus[data_w*3 +:data_w];
assign c20ibus[temp_w*4 +:temp_w] = v1179obus[temp_w*0 +:temp_w];
assign v1179ibus[data_w*0 +:data_w] = c20obus[data_w*4 +:data_w];
assign c20ibus[temp_w*5 +:temp_w] = v1268obus[temp_w*0 +:temp_w];
assign v1268ibus[data_w*0 +:data_w] = c20obus[data_w*5 +:data_w];
assign c21ibus[temp_w*0 +:temp_w] = v115obus[temp_w*0 +:temp_w];
assign v115ibus[data_w*0 +:data_w] = c21obus[data_w*0 +:data_w];
assign c21ibus[temp_w*1 +:temp_w] = v286obus[temp_w*0 +:temp_w];
assign v286ibus[data_w*0 +:data_w] = c21obus[data_w*1 +:data_w];
assign c21ibus[temp_w*2 +:temp_w] = v844obus[temp_w*0 +:temp_w];
assign v844ibus[data_w*0 +:data_w] = c21obus[data_w*2 +:data_w];
assign c21ibus[temp_w*3 +:temp_w] = v872obus[temp_w*0 +:temp_w];
assign v872ibus[data_w*0 +:data_w] = c21obus[data_w*3 +:data_w];
assign c21ibus[temp_w*4 +:temp_w] = v1180obus[temp_w*0 +:temp_w];
assign v1180ibus[data_w*0 +:data_w] = c21obus[data_w*4 +:data_w];
assign c21ibus[temp_w*5 +:temp_w] = v1269obus[temp_w*0 +:temp_w];
assign v1269ibus[data_w*0 +:data_w] = c21obus[data_w*5 +:data_w];
assign c22ibus[temp_w*0 +:temp_w] = v116obus[temp_w*0 +:temp_w];
assign v116ibus[data_w*0 +:data_w] = c22obus[data_w*0 +:data_w];
assign c22ibus[temp_w*1 +:temp_w] = v287obus[temp_w*0 +:temp_w];
assign v287ibus[data_w*0 +:data_w] = c22obus[data_w*1 +:data_w];
assign c22ibus[temp_w*2 +:temp_w] = v845obus[temp_w*0 +:temp_w];
assign v845ibus[data_w*0 +:data_w] = c22obus[data_w*2 +:data_w];
assign c22ibus[temp_w*3 +:temp_w] = v873obus[temp_w*0 +:temp_w];
assign v873ibus[data_w*0 +:data_w] = c22obus[data_w*3 +:data_w];
assign c22ibus[temp_w*4 +:temp_w] = v1181obus[temp_w*0 +:temp_w];
assign v1181ibus[data_w*0 +:data_w] = c22obus[data_w*4 +:data_w];
assign c22ibus[temp_w*5 +:temp_w] = v1270obus[temp_w*0 +:temp_w];
assign v1270ibus[data_w*0 +:data_w] = c22obus[data_w*5 +:data_w];
assign c23ibus[temp_w*0 +:temp_w] = v117obus[temp_w*0 +:temp_w];
assign v117ibus[data_w*0 +:data_w] = c23obus[data_w*0 +:data_w];
assign c23ibus[temp_w*1 +:temp_w] = v192obus[temp_w*0 +:temp_w];
assign v192ibus[data_w*0 +:data_w] = c23obus[data_w*1 +:data_w];
assign c23ibus[temp_w*2 +:temp_w] = v846obus[temp_w*0 +:temp_w];
assign v846ibus[data_w*0 +:data_w] = c23obus[data_w*2 +:data_w];
assign c23ibus[temp_w*3 +:temp_w] = v874obus[temp_w*0 +:temp_w];
assign v874ibus[data_w*0 +:data_w] = c23obus[data_w*3 +:data_w];
assign c23ibus[temp_w*4 +:temp_w] = v1182obus[temp_w*0 +:temp_w];
assign v1182ibus[data_w*0 +:data_w] = c23obus[data_w*4 +:data_w];
assign c23ibus[temp_w*5 +:temp_w] = v1271obus[temp_w*0 +:temp_w];
assign v1271ibus[data_w*0 +:data_w] = c23obus[data_w*5 +:data_w];
assign c24ibus[temp_w*0 +:temp_w] = v118obus[temp_w*0 +:temp_w];
assign v118ibus[data_w*0 +:data_w] = c24obus[data_w*0 +:data_w];
assign c24ibus[temp_w*1 +:temp_w] = v193obus[temp_w*0 +:temp_w];
assign v193ibus[data_w*0 +:data_w] = c24obus[data_w*1 +:data_w];
assign c24ibus[temp_w*2 +:temp_w] = v847obus[temp_w*0 +:temp_w];
assign v847ibus[data_w*0 +:data_w] = c24obus[data_w*2 +:data_w];
assign c24ibus[temp_w*3 +:temp_w] = v875obus[temp_w*0 +:temp_w];
assign v875ibus[data_w*0 +:data_w] = c24obus[data_w*3 +:data_w];
assign c24ibus[temp_w*4 +:temp_w] = v1183obus[temp_w*0 +:temp_w];
assign v1183ibus[data_w*0 +:data_w] = c24obus[data_w*4 +:data_w];
assign c24ibus[temp_w*5 +:temp_w] = v1272obus[temp_w*0 +:temp_w];
assign v1272ibus[data_w*0 +:data_w] = c24obus[data_w*5 +:data_w];
assign c25ibus[temp_w*0 +:temp_w] = v119obus[temp_w*0 +:temp_w];
assign v119ibus[data_w*0 +:data_w] = c25obus[data_w*0 +:data_w];
assign c25ibus[temp_w*1 +:temp_w] = v194obus[temp_w*0 +:temp_w];
assign v194ibus[data_w*0 +:data_w] = c25obus[data_w*1 +:data_w];
assign c25ibus[temp_w*2 +:temp_w] = v848obus[temp_w*0 +:temp_w];
assign v848ibus[data_w*0 +:data_w] = c25obus[data_w*2 +:data_w];
assign c25ibus[temp_w*3 +:temp_w] = v876obus[temp_w*0 +:temp_w];
assign v876ibus[data_w*0 +:data_w] = c25obus[data_w*3 +:data_w];
assign c25ibus[temp_w*4 +:temp_w] = v1184obus[temp_w*0 +:temp_w];
assign v1184ibus[data_w*0 +:data_w] = c25obus[data_w*4 +:data_w];
assign c25ibus[temp_w*5 +:temp_w] = v1273obus[temp_w*0 +:temp_w];
assign v1273ibus[data_w*0 +:data_w] = c25obus[data_w*5 +:data_w];
assign c26ibus[temp_w*0 +:temp_w] = v120obus[temp_w*0 +:temp_w];
assign v120ibus[data_w*0 +:data_w] = c26obus[data_w*0 +:data_w];
assign c26ibus[temp_w*1 +:temp_w] = v195obus[temp_w*0 +:temp_w];
assign v195ibus[data_w*0 +:data_w] = c26obus[data_w*1 +:data_w];
assign c26ibus[temp_w*2 +:temp_w] = v849obus[temp_w*0 +:temp_w];
assign v849ibus[data_w*0 +:data_w] = c26obus[data_w*2 +:data_w];
assign c26ibus[temp_w*3 +:temp_w] = v877obus[temp_w*0 +:temp_w];
assign v877ibus[data_w*0 +:data_w] = c26obus[data_w*3 +:data_w];
assign c26ibus[temp_w*4 +:temp_w] = v1185obus[temp_w*0 +:temp_w];
assign v1185ibus[data_w*0 +:data_w] = c26obus[data_w*4 +:data_w];
assign c26ibus[temp_w*5 +:temp_w] = v1274obus[temp_w*0 +:temp_w];
assign v1274ibus[data_w*0 +:data_w] = c26obus[data_w*5 +:data_w];
assign c27ibus[temp_w*0 +:temp_w] = v121obus[temp_w*0 +:temp_w];
assign v121ibus[data_w*0 +:data_w] = c27obus[data_w*0 +:data_w];
assign c27ibus[temp_w*1 +:temp_w] = v196obus[temp_w*0 +:temp_w];
assign v196ibus[data_w*0 +:data_w] = c27obus[data_w*1 +:data_w];
assign c27ibus[temp_w*2 +:temp_w] = v850obus[temp_w*0 +:temp_w];
assign v850ibus[data_w*0 +:data_w] = c27obus[data_w*2 +:data_w];
assign c27ibus[temp_w*3 +:temp_w] = v878obus[temp_w*0 +:temp_w];
assign v878ibus[data_w*0 +:data_w] = c27obus[data_w*3 +:data_w];
assign c27ibus[temp_w*4 +:temp_w] = v1186obus[temp_w*0 +:temp_w];
assign v1186ibus[data_w*0 +:data_w] = c27obus[data_w*4 +:data_w];
assign c27ibus[temp_w*5 +:temp_w] = v1275obus[temp_w*0 +:temp_w];
assign v1275ibus[data_w*0 +:data_w] = c27obus[data_w*5 +:data_w];
assign c28ibus[temp_w*0 +:temp_w] = v122obus[temp_w*0 +:temp_w];
assign v122ibus[data_w*0 +:data_w] = c28obus[data_w*0 +:data_w];
assign c28ibus[temp_w*1 +:temp_w] = v197obus[temp_w*0 +:temp_w];
assign v197ibus[data_w*0 +:data_w] = c28obus[data_w*1 +:data_w];
assign c28ibus[temp_w*2 +:temp_w] = v851obus[temp_w*0 +:temp_w];
assign v851ibus[data_w*0 +:data_w] = c28obus[data_w*2 +:data_w];
assign c28ibus[temp_w*3 +:temp_w] = v879obus[temp_w*0 +:temp_w];
assign v879ibus[data_w*0 +:data_w] = c28obus[data_w*3 +:data_w];
assign c28ibus[temp_w*4 +:temp_w] = v1187obus[temp_w*0 +:temp_w];
assign v1187ibus[data_w*0 +:data_w] = c28obus[data_w*4 +:data_w];
assign c28ibus[temp_w*5 +:temp_w] = v1276obus[temp_w*0 +:temp_w];
assign v1276ibus[data_w*0 +:data_w] = c28obus[data_w*5 +:data_w];
assign c29ibus[temp_w*0 +:temp_w] = v123obus[temp_w*0 +:temp_w];
assign v123ibus[data_w*0 +:data_w] = c29obus[data_w*0 +:data_w];
assign c29ibus[temp_w*1 +:temp_w] = v198obus[temp_w*0 +:temp_w];
assign v198ibus[data_w*0 +:data_w] = c29obus[data_w*1 +:data_w];
assign c29ibus[temp_w*2 +:temp_w] = v852obus[temp_w*0 +:temp_w];
assign v852ibus[data_w*0 +:data_w] = c29obus[data_w*2 +:data_w];
assign c29ibus[temp_w*3 +:temp_w] = v880obus[temp_w*0 +:temp_w];
assign v880ibus[data_w*0 +:data_w] = c29obus[data_w*3 +:data_w];
assign c29ibus[temp_w*4 +:temp_w] = v1188obus[temp_w*0 +:temp_w];
assign v1188ibus[data_w*0 +:data_w] = c29obus[data_w*4 +:data_w];
assign c29ibus[temp_w*5 +:temp_w] = v1277obus[temp_w*0 +:temp_w];
assign v1277ibus[data_w*0 +:data_w] = c29obus[data_w*5 +:data_w];
assign c30ibus[temp_w*0 +:temp_w] = v124obus[temp_w*0 +:temp_w];
assign v124ibus[data_w*0 +:data_w] = c30obus[data_w*0 +:data_w];
assign c30ibus[temp_w*1 +:temp_w] = v199obus[temp_w*0 +:temp_w];
assign v199ibus[data_w*0 +:data_w] = c30obus[data_w*1 +:data_w];
assign c30ibus[temp_w*2 +:temp_w] = v853obus[temp_w*0 +:temp_w];
assign v853ibus[data_w*0 +:data_w] = c30obus[data_w*2 +:data_w];
assign c30ibus[temp_w*3 +:temp_w] = v881obus[temp_w*0 +:temp_w];
assign v881ibus[data_w*0 +:data_w] = c30obus[data_w*3 +:data_w];
assign c30ibus[temp_w*4 +:temp_w] = v1189obus[temp_w*0 +:temp_w];
assign v1189ibus[data_w*0 +:data_w] = c30obus[data_w*4 +:data_w];
assign c30ibus[temp_w*5 +:temp_w] = v1278obus[temp_w*0 +:temp_w];
assign v1278ibus[data_w*0 +:data_w] = c30obus[data_w*5 +:data_w];
assign c31ibus[temp_w*0 +:temp_w] = v125obus[temp_w*0 +:temp_w];
assign v125ibus[data_w*0 +:data_w] = c31obus[data_w*0 +:data_w];
assign c31ibus[temp_w*1 +:temp_w] = v200obus[temp_w*0 +:temp_w];
assign v200ibus[data_w*0 +:data_w] = c31obus[data_w*1 +:data_w];
assign c31ibus[temp_w*2 +:temp_w] = v854obus[temp_w*0 +:temp_w];
assign v854ibus[data_w*0 +:data_w] = c31obus[data_w*2 +:data_w];
assign c31ibus[temp_w*3 +:temp_w] = v882obus[temp_w*0 +:temp_w];
assign v882ibus[data_w*0 +:data_w] = c31obus[data_w*3 +:data_w];
assign c31ibus[temp_w*4 +:temp_w] = v1190obus[temp_w*0 +:temp_w];
assign v1190ibus[data_w*0 +:data_w] = c31obus[data_w*4 +:data_w];
assign c31ibus[temp_w*5 +:temp_w] = v1279obus[temp_w*0 +:temp_w];
assign v1279ibus[data_w*0 +:data_w] = c31obus[data_w*5 +:data_w];
assign c32ibus[temp_w*0 +:temp_w] = v126obus[temp_w*0 +:temp_w];
assign v126ibus[data_w*0 +:data_w] = c32obus[data_w*0 +:data_w];
assign c32ibus[temp_w*1 +:temp_w] = v201obus[temp_w*0 +:temp_w];
assign v201ibus[data_w*0 +:data_w] = c32obus[data_w*1 +:data_w];
assign c32ibus[temp_w*2 +:temp_w] = v855obus[temp_w*0 +:temp_w];
assign v855ibus[data_w*0 +:data_w] = c32obus[data_w*2 +:data_w];
assign c32ibus[temp_w*3 +:temp_w] = v883obus[temp_w*0 +:temp_w];
assign v883ibus[data_w*0 +:data_w] = c32obus[data_w*3 +:data_w];
assign c32ibus[temp_w*4 +:temp_w] = v1191obus[temp_w*0 +:temp_w];
assign v1191ibus[data_w*0 +:data_w] = c32obus[data_w*4 +:data_w];
assign c32ibus[temp_w*5 +:temp_w] = v1280obus[temp_w*0 +:temp_w];
assign v1280ibus[data_w*0 +:data_w] = c32obus[data_w*5 +:data_w];
assign c33ibus[temp_w*0 +:temp_w] = v127obus[temp_w*0 +:temp_w];
assign v127ibus[data_w*0 +:data_w] = c33obus[data_w*0 +:data_w];
assign c33ibus[temp_w*1 +:temp_w] = v202obus[temp_w*0 +:temp_w];
assign v202ibus[data_w*0 +:data_w] = c33obus[data_w*1 +:data_w];
assign c33ibus[temp_w*2 +:temp_w] = v856obus[temp_w*0 +:temp_w];
assign v856ibus[data_w*0 +:data_w] = c33obus[data_w*2 +:data_w];
assign c33ibus[temp_w*3 +:temp_w] = v884obus[temp_w*0 +:temp_w];
assign v884ibus[data_w*0 +:data_w] = c33obus[data_w*3 +:data_w];
assign c33ibus[temp_w*4 +:temp_w] = v1192obus[temp_w*0 +:temp_w];
assign v1192ibus[data_w*0 +:data_w] = c33obus[data_w*4 +:data_w];
assign c33ibus[temp_w*5 +:temp_w] = v1281obus[temp_w*0 +:temp_w];
assign v1281ibus[data_w*0 +:data_w] = c33obus[data_w*5 +:data_w];
assign c34ibus[temp_w*0 +:temp_w] = v128obus[temp_w*0 +:temp_w];
assign v128ibus[data_w*0 +:data_w] = c34obus[data_w*0 +:data_w];
assign c34ibus[temp_w*1 +:temp_w] = v203obus[temp_w*0 +:temp_w];
assign v203ibus[data_w*0 +:data_w] = c34obus[data_w*1 +:data_w];
assign c34ibus[temp_w*2 +:temp_w] = v857obus[temp_w*0 +:temp_w];
assign v857ibus[data_w*0 +:data_w] = c34obus[data_w*2 +:data_w];
assign c34ibus[temp_w*3 +:temp_w] = v885obus[temp_w*0 +:temp_w];
assign v885ibus[data_w*0 +:data_w] = c34obus[data_w*3 +:data_w];
assign c34ibus[temp_w*4 +:temp_w] = v1193obus[temp_w*0 +:temp_w];
assign v1193ibus[data_w*0 +:data_w] = c34obus[data_w*4 +:data_w];
assign c34ibus[temp_w*5 +:temp_w] = v1282obus[temp_w*0 +:temp_w];
assign v1282ibus[data_w*0 +:data_w] = c34obus[data_w*5 +:data_w];
assign c35ibus[temp_w*0 +:temp_w] = v129obus[temp_w*0 +:temp_w];
assign v129ibus[data_w*0 +:data_w] = c35obus[data_w*0 +:data_w];
assign c35ibus[temp_w*1 +:temp_w] = v204obus[temp_w*0 +:temp_w];
assign v204ibus[data_w*0 +:data_w] = c35obus[data_w*1 +:data_w];
assign c35ibus[temp_w*2 +:temp_w] = v858obus[temp_w*0 +:temp_w];
assign v858ibus[data_w*0 +:data_w] = c35obus[data_w*2 +:data_w];
assign c35ibus[temp_w*3 +:temp_w] = v886obus[temp_w*0 +:temp_w];
assign v886ibus[data_w*0 +:data_w] = c35obus[data_w*3 +:data_w];
assign c35ibus[temp_w*4 +:temp_w] = v1194obus[temp_w*0 +:temp_w];
assign v1194ibus[data_w*0 +:data_w] = c35obus[data_w*4 +:data_w];
assign c35ibus[temp_w*5 +:temp_w] = v1283obus[temp_w*0 +:temp_w];
assign v1283ibus[data_w*0 +:data_w] = c35obus[data_w*5 +:data_w];
assign c36ibus[temp_w*0 +:temp_w] = v130obus[temp_w*0 +:temp_w];
assign v130ibus[data_w*0 +:data_w] = c36obus[data_w*0 +:data_w];
assign c36ibus[temp_w*1 +:temp_w] = v205obus[temp_w*0 +:temp_w];
assign v205ibus[data_w*0 +:data_w] = c36obus[data_w*1 +:data_w];
assign c36ibus[temp_w*2 +:temp_w] = v859obus[temp_w*0 +:temp_w];
assign v859ibus[data_w*0 +:data_w] = c36obus[data_w*2 +:data_w];
assign c36ibus[temp_w*3 +:temp_w] = v887obus[temp_w*0 +:temp_w];
assign v887ibus[data_w*0 +:data_w] = c36obus[data_w*3 +:data_w];
assign c36ibus[temp_w*4 +:temp_w] = v1195obus[temp_w*0 +:temp_w];
assign v1195ibus[data_w*0 +:data_w] = c36obus[data_w*4 +:data_w];
assign c36ibus[temp_w*5 +:temp_w] = v1284obus[temp_w*0 +:temp_w];
assign v1284ibus[data_w*0 +:data_w] = c36obus[data_w*5 +:data_w];
assign c37ibus[temp_w*0 +:temp_w] = v131obus[temp_w*0 +:temp_w];
assign v131ibus[data_w*0 +:data_w] = c37obus[data_w*0 +:data_w];
assign c37ibus[temp_w*1 +:temp_w] = v206obus[temp_w*0 +:temp_w];
assign v206ibus[data_w*0 +:data_w] = c37obus[data_w*1 +:data_w];
assign c37ibus[temp_w*2 +:temp_w] = v860obus[temp_w*0 +:temp_w];
assign v860ibus[data_w*0 +:data_w] = c37obus[data_w*2 +:data_w];
assign c37ibus[temp_w*3 +:temp_w] = v888obus[temp_w*0 +:temp_w];
assign v888ibus[data_w*0 +:data_w] = c37obus[data_w*3 +:data_w];
assign c37ibus[temp_w*4 +:temp_w] = v1196obus[temp_w*0 +:temp_w];
assign v1196ibus[data_w*0 +:data_w] = c37obus[data_w*4 +:data_w];
assign c37ibus[temp_w*5 +:temp_w] = v1285obus[temp_w*0 +:temp_w];
assign v1285ibus[data_w*0 +:data_w] = c37obus[data_w*5 +:data_w];
assign c38ibus[temp_w*0 +:temp_w] = v132obus[temp_w*0 +:temp_w];
assign v132ibus[data_w*0 +:data_w] = c38obus[data_w*0 +:data_w];
assign c38ibus[temp_w*1 +:temp_w] = v207obus[temp_w*0 +:temp_w];
assign v207ibus[data_w*0 +:data_w] = c38obus[data_w*1 +:data_w];
assign c38ibus[temp_w*2 +:temp_w] = v861obus[temp_w*0 +:temp_w];
assign v861ibus[data_w*0 +:data_w] = c38obus[data_w*2 +:data_w];
assign c38ibus[temp_w*3 +:temp_w] = v889obus[temp_w*0 +:temp_w];
assign v889ibus[data_w*0 +:data_w] = c38obus[data_w*3 +:data_w];
assign c38ibus[temp_w*4 +:temp_w] = v1197obus[temp_w*0 +:temp_w];
assign v1197ibus[data_w*0 +:data_w] = c38obus[data_w*4 +:data_w];
assign c38ibus[temp_w*5 +:temp_w] = v1286obus[temp_w*0 +:temp_w];
assign v1286ibus[data_w*0 +:data_w] = c38obus[data_w*5 +:data_w];
assign c39ibus[temp_w*0 +:temp_w] = v133obus[temp_w*0 +:temp_w];
assign v133ibus[data_w*0 +:data_w] = c39obus[data_w*0 +:data_w];
assign c39ibus[temp_w*1 +:temp_w] = v208obus[temp_w*0 +:temp_w];
assign v208ibus[data_w*0 +:data_w] = c39obus[data_w*1 +:data_w];
assign c39ibus[temp_w*2 +:temp_w] = v862obus[temp_w*0 +:temp_w];
assign v862ibus[data_w*0 +:data_w] = c39obus[data_w*2 +:data_w];
assign c39ibus[temp_w*3 +:temp_w] = v890obus[temp_w*0 +:temp_w];
assign v890ibus[data_w*0 +:data_w] = c39obus[data_w*3 +:data_w];
assign c39ibus[temp_w*4 +:temp_w] = v1198obus[temp_w*0 +:temp_w];
assign v1198ibus[data_w*0 +:data_w] = c39obus[data_w*4 +:data_w];
assign c39ibus[temp_w*5 +:temp_w] = v1287obus[temp_w*0 +:temp_w];
assign v1287ibus[data_w*0 +:data_w] = c39obus[data_w*5 +:data_w];
assign c40ibus[temp_w*0 +:temp_w] = v134obus[temp_w*0 +:temp_w];
assign v134ibus[data_w*0 +:data_w] = c40obus[data_w*0 +:data_w];
assign c40ibus[temp_w*1 +:temp_w] = v209obus[temp_w*0 +:temp_w];
assign v209ibus[data_w*0 +:data_w] = c40obus[data_w*1 +:data_w];
assign c40ibus[temp_w*2 +:temp_w] = v863obus[temp_w*0 +:temp_w];
assign v863ibus[data_w*0 +:data_w] = c40obus[data_w*2 +:data_w];
assign c40ibus[temp_w*3 +:temp_w] = v891obus[temp_w*0 +:temp_w];
assign v891ibus[data_w*0 +:data_w] = c40obus[data_w*3 +:data_w];
assign c40ibus[temp_w*4 +:temp_w] = v1199obus[temp_w*0 +:temp_w];
assign v1199ibus[data_w*0 +:data_w] = c40obus[data_w*4 +:data_w];
assign c40ibus[temp_w*5 +:temp_w] = v1288obus[temp_w*0 +:temp_w];
assign v1288ibus[data_w*0 +:data_w] = c40obus[data_w*5 +:data_w];
assign c41ibus[temp_w*0 +:temp_w] = v135obus[temp_w*0 +:temp_w];
assign v135ibus[data_w*0 +:data_w] = c41obus[data_w*0 +:data_w];
assign c41ibus[temp_w*1 +:temp_w] = v210obus[temp_w*0 +:temp_w];
assign v210ibus[data_w*0 +:data_w] = c41obus[data_w*1 +:data_w];
assign c41ibus[temp_w*2 +:temp_w] = v768obus[temp_w*0 +:temp_w];
assign v768ibus[data_w*0 +:data_w] = c41obus[data_w*2 +:data_w];
assign c41ibus[temp_w*3 +:temp_w] = v892obus[temp_w*0 +:temp_w];
assign v892ibus[data_w*0 +:data_w] = c41obus[data_w*3 +:data_w];
assign c41ibus[temp_w*4 +:temp_w] = v1200obus[temp_w*0 +:temp_w];
assign v1200ibus[data_w*0 +:data_w] = c41obus[data_w*4 +:data_w];
assign c41ibus[temp_w*5 +:temp_w] = v1289obus[temp_w*0 +:temp_w];
assign v1289ibus[data_w*0 +:data_w] = c41obus[data_w*5 +:data_w];
assign c42ibus[temp_w*0 +:temp_w] = v136obus[temp_w*0 +:temp_w];
assign v136ibus[data_w*0 +:data_w] = c42obus[data_w*0 +:data_w];
assign c42ibus[temp_w*1 +:temp_w] = v211obus[temp_w*0 +:temp_w];
assign v211ibus[data_w*0 +:data_w] = c42obus[data_w*1 +:data_w];
assign c42ibus[temp_w*2 +:temp_w] = v769obus[temp_w*0 +:temp_w];
assign v769ibus[data_w*0 +:data_w] = c42obus[data_w*2 +:data_w];
assign c42ibus[temp_w*3 +:temp_w] = v893obus[temp_w*0 +:temp_w];
assign v893ibus[data_w*0 +:data_w] = c42obus[data_w*3 +:data_w];
assign c42ibus[temp_w*4 +:temp_w] = v1201obus[temp_w*0 +:temp_w];
assign v1201ibus[data_w*0 +:data_w] = c42obus[data_w*4 +:data_w];
assign c42ibus[temp_w*5 +:temp_w] = v1290obus[temp_w*0 +:temp_w];
assign v1290ibus[data_w*0 +:data_w] = c42obus[data_w*5 +:data_w];
assign c43ibus[temp_w*0 +:temp_w] = v137obus[temp_w*0 +:temp_w];
assign v137ibus[data_w*0 +:data_w] = c43obus[data_w*0 +:data_w];
assign c43ibus[temp_w*1 +:temp_w] = v212obus[temp_w*0 +:temp_w];
assign v212ibus[data_w*0 +:data_w] = c43obus[data_w*1 +:data_w];
assign c43ibus[temp_w*2 +:temp_w] = v770obus[temp_w*0 +:temp_w];
assign v770ibus[data_w*0 +:data_w] = c43obus[data_w*2 +:data_w];
assign c43ibus[temp_w*3 +:temp_w] = v894obus[temp_w*0 +:temp_w];
assign v894ibus[data_w*0 +:data_w] = c43obus[data_w*3 +:data_w];
assign c43ibus[temp_w*4 +:temp_w] = v1202obus[temp_w*0 +:temp_w];
assign v1202ibus[data_w*0 +:data_w] = c43obus[data_w*4 +:data_w];
assign c43ibus[temp_w*5 +:temp_w] = v1291obus[temp_w*0 +:temp_w];
assign v1291ibus[data_w*0 +:data_w] = c43obus[data_w*5 +:data_w];
assign c44ibus[temp_w*0 +:temp_w] = v138obus[temp_w*0 +:temp_w];
assign v138ibus[data_w*0 +:data_w] = c44obus[data_w*0 +:data_w];
assign c44ibus[temp_w*1 +:temp_w] = v213obus[temp_w*0 +:temp_w];
assign v213ibus[data_w*0 +:data_w] = c44obus[data_w*1 +:data_w];
assign c44ibus[temp_w*2 +:temp_w] = v771obus[temp_w*0 +:temp_w];
assign v771ibus[data_w*0 +:data_w] = c44obus[data_w*2 +:data_w];
assign c44ibus[temp_w*3 +:temp_w] = v895obus[temp_w*0 +:temp_w];
assign v895ibus[data_w*0 +:data_w] = c44obus[data_w*3 +:data_w];
assign c44ibus[temp_w*4 +:temp_w] = v1203obus[temp_w*0 +:temp_w];
assign v1203ibus[data_w*0 +:data_w] = c44obus[data_w*4 +:data_w];
assign c44ibus[temp_w*5 +:temp_w] = v1292obus[temp_w*0 +:temp_w];
assign v1292ibus[data_w*0 +:data_w] = c44obus[data_w*5 +:data_w];
assign c45ibus[temp_w*0 +:temp_w] = v139obus[temp_w*0 +:temp_w];
assign v139ibus[data_w*0 +:data_w] = c45obus[data_w*0 +:data_w];
assign c45ibus[temp_w*1 +:temp_w] = v214obus[temp_w*0 +:temp_w];
assign v214ibus[data_w*0 +:data_w] = c45obus[data_w*1 +:data_w];
assign c45ibus[temp_w*2 +:temp_w] = v772obus[temp_w*0 +:temp_w];
assign v772ibus[data_w*0 +:data_w] = c45obus[data_w*2 +:data_w];
assign c45ibus[temp_w*3 +:temp_w] = v896obus[temp_w*0 +:temp_w];
assign v896ibus[data_w*0 +:data_w] = c45obus[data_w*3 +:data_w];
assign c45ibus[temp_w*4 +:temp_w] = v1204obus[temp_w*0 +:temp_w];
assign v1204ibus[data_w*0 +:data_w] = c45obus[data_w*4 +:data_w];
assign c45ibus[temp_w*5 +:temp_w] = v1293obus[temp_w*0 +:temp_w];
assign v1293ibus[data_w*0 +:data_w] = c45obus[data_w*5 +:data_w];
assign c46ibus[temp_w*0 +:temp_w] = v140obus[temp_w*0 +:temp_w];
assign v140ibus[data_w*0 +:data_w] = c46obus[data_w*0 +:data_w];
assign c46ibus[temp_w*1 +:temp_w] = v215obus[temp_w*0 +:temp_w];
assign v215ibus[data_w*0 +:data_w] = c46obus[data_w*1 +:data_w];
assign c46ibus[temp_w*2 +:temp_w] = v773obus[temp_w*0 +:temp_w];
assign v773ibus[data_w*0 +:data_w] = c46obus[data_w*2 +:data_w];
assign c46ibus[temp_w*3 +:temp_w] = v897obus[temp_w*0 +:temp_w];
assign v897ibus[data_w*0 +:data_w] = c46obus[data_w*3 +:data_w];
assign c46ibus[temp_w*4 +:temp_w] = v1205obus[temp_w*0 +:temp_w];
assign v1205ibus[data_w*0 +:data_w] = c46obus[data_w*4 +:data_w];
assign c46ibus[temp_w*5 +:temp_w] = v1294obus[temp_w*0 +:temp_w];
assign v1294ibus[data_w*0 +:data_w] = c46obus[data_w*5 +:data_w];
assign c47ibus[temp_w*0 +:temp_w] = v141obus[temp_w*0 +:temp_w];
assign v141ibus[data_w*0 +:data_w] = c47obus[data_w*0 +:data_w];
assign c47ibus[temp_w*1 +:temp_w] = v216obus[temp_w*0 +:temp_w];
assign v216ibus[data_w*0 +:data_w] = c47obus[data_w*1 +:data_w];
assign c47ibus[temp_w*2 +:temp_w] = v774obus[temp_w*0 +:temp_w];
assign v774ibus[data_w*0 +:data_w] = c47obus[data_w*2 +:data_w];
assign c47ibus[temp_w*3 +:temp_w] = v898obus[temp_w*0 +:temp_w];
assign v898ibus[data_w*0 +:data_w] = c47obus[data_w*3 +:data_w];
assign c47ibus[temp_w*4 +:temp_w] = v1206obus[temp_w*0 +:temp_w];
assign v1206ibus[data_w*0 +:data_w] = c47obus[data_w*4 +:data_w];
assign c47ibus[temp_w*5 +:temp_w] = v1295obus[temp_w*0 +:temp_w];
assign v1295ibus[data_w*0 +:data_w] = c47obus[data_w*5 +:data_w];
assign c48ibus[temp_w*0 +:temp_w] = v142obus[temp_w*0 +:temp_w];
assign v142ibus[data_w*0 +:data_w] = c48obus[data_w*0 +:data_w];
assign c48ibus[temp_w*1 +:temp_w] = v217obus[temp_w*0 +:temp_w];
assign v217ibus[data_w*0 +:data_w] = c48obus[data_w*1 +:data_w];
assign c48ibus[temp_w*2 +:temp_w] = v775obus[temp_w*0 +:temp_w];
assign v775ibus[data_w*0 +:data_w] = c48obus[data_w*2 +:data_w];
assign c48ibus[temp_w*3 +:temp_w] = v899obus[temp_w*0 +:temp_w];
assign v899ibus[data_w*0 +:data_w] = c48obus[data_w*3 +:data_w];
assign c48ibus[temp_w*4 +:temp_w] = v1207obus[temp_w*0 +:temp_w];
assign v1207ibus[data_w*0 +:data_w] = c48obus[data_w*4 +:data_w];
assign c48ibus[temp_w*5 +:temp_w] = v1296obus[temp_w*0 +:temp_w];
assign v1296ibus[data_w*0 +:data_w] = c48obus[data_w*5 +:data_w];
assign c49ibus[temp_w*0 +:temp_w] = v143obus[temp_w*0 +:temp_w];
assign v143ibus[data_w*0 +:data_w] = c49obus[data_w*0 +:data_w];
assign c49ibus[temp_w*1 +:temp_w] = v218obus[temp_w*0 +:temp_w];
assign v218ibus[data_w*0 +:data_w] = c49obus[data_w*1 +:data_w];
assign c49ibus[temp_w*2 +:temp_w] = v776obus[temp_w*0 +:temp_w];
assign v776ibus[data_w*0 +:data_w] = c49obus[data_w*2 +:data_w];
assign c49ibus[temp_w*3 +:temp_w] = v900obus[temp_w*0 +:temp_w];
assign v900ibus[data_w*0 +:data_w] = c49obus[data_w*3 +:data_w];
assign c49ibus[temp_w*4 +:temp_w] = v1208obus[temp_w*0 +:temp_w];
assign v1208ibus[data_w*0 +:data_w] = c49obus[data_w*4 +:data_w];
assign c49ibus[temp_w*5 +:temp_w] = v1297obus[temp_w*0 +:temp_w];
assign v1297ibus[data_w*0 +:data_w] = c49obus[data_w*5 +:data_w];
assign c50ibus[temp_w*0 +:temp_w] = v144obus[temp_w*0 +:temp_w];
assign v144ibus[data_w*0 +:data_w] = c50obus[data_w*0 +:data_w];
assign c50ibus[temp_w*1 +:temp_w] = v219obus[temp_w*0 +:temp_w];
assign v219ibus[data_w*0 +:data_w] = c50obus[data_w*1 +:data_w];
assign c50ibus[temp_w*2 +:temp_w] = v777obus[temp_w*0 +:temp_w];
assign v777ibus[data_w*0 +:data_w] = c50obus[data_w*2 +:data_w];
assign c50ibus[temp_w*3 +:temp_w] = v901obus[temp_w*0 +:temp_w];
assign v901ibus[data_w*0 +:data_w] = c50obus[data_w*3 +:data_w];
assign c50ibus[temp_w*4 +:temp_w] = v1209obus[temp_w*0 +:temp_w];
assign v1209ibus[data_w*0 +:data_w] = c50obus[data_w*4 +:data_w];
assign c50ibus[temp_w*5 +:temp_w] = v1298obus[temp_w*0 +:temp_w];
assign v1298ibus[data_w*0 +:data_w] = c50obus[data_w*5 +:data_w];
assign c51ibus[temp_w*0 +:temp_w] = v145obus[temp_w*0 +:temp_w];
assign v145ibus[data_w*0 +:data_w] = c51obus[data_w*0 +:data_w];
assign c51ibus[temp_w*1 +:temp_w] = v220obus[temp_w*0 +:temp_w];
assign v220ibus[data_w*0 +:data_w] = c51obus[data_w*1 +:data_w];
assign c51ibus[temp_w*2 +:temp_w] = v778obus[temp_w*0 +:temp_w];
assign v778ibus[data_w*0 +:data_w] = c51obus[data_w*2 +:data_w];
assign c51ibus[temp_w*3 +:temp_w] = v902obus[temp_w*0 +:temp_w];
assign v902ibus[data_w*0 +:data_w] = c51obus[data_w*3 +:data_w];
assign c51ibus[temp_w*4 +:temp_w] = v1210obus[temp_w*0 +:temp_w];
assign v1210ibus[data_w*0 +:data_w] = c51obus[data_w*4 +:data_w];
assign c51ibus[temp_w*5 +:temp_w] = v1299obus[temp_w*0 +:temp_w];
assign v1299ibus[data_w*0 +:data_w] = c51obus[data_w*5 +:data_w];
assign c52ibus[temp_w*0 +:temp_w] = v146obus[temp_w*0 +:temp_w];
assign v146ibus[data_w*0 +:data_w] = c52obus[data_w*0 +:data_w];
assign c52ibus[temp_w*1 +:temp_w] = v221obus[temp_w*0 +:temp_w];
assign v221ibus[data_w*0 +:data_w] = c52obus[data_w*1 +:data_w];
assign c52ibus[temp_w*2 +:temp_w] = v779obus[temp_w*0 +:temp_w];
assign v779ibus[data_w*0 +:data_w] = c52obus[data_w*2 +:data_w];
assign c52ibus[temp_w*3 +:temp_w] = v903obus[temp_w*0 +:temp_w];
assign v903ibus[data_w*0 +:data_w] = c52obus[data_w*3 +:data_w];
assign c52ibus[temp_w*4 +:temp_w] = v1211obus[temp_w*0 +:temp_w];
assign v1211ibus[data_w*0 +:data_w] = c52obus[data_w*4 +:data_w];
assign c52ibus[temp_w*5 +:temp_w] = v1300obus[temp_w*0 +:temp_w];
assign v1300ibus[data_w*0 +:data_w] = c52obus[data_w*5 +:data_w];
assign c53ibus[temp_w*0 +:temp_w] = v147obus[temp_w*0 +:temp_w];
assign v147ibus[data_w*0 +:data_w] = c53obus[data_w*0 +:data_w];
assign c53ibus[temp_w*1 +:temp_w] = v222obus[temp_w*0 +:temp_w];
assign v222ibus[data_w*0 +:data_w] = c53obus[data_w*1 +:data_w];
assign c53ibus[temp_w*2 +:temp_w] = v780obus[temp_w*0 +:temp_w];
assign v780ibus[data_w*0 +:data_w] = c53obus[data_w*2 +:data_w];
assign c53ibus[temp_w*3 +:temp_w] = v904obus[temp_w*0 +:temp_w];
assign v904ibus[data_w*0 +:data_w] = c53obus[data_w*3 +:data_w];
assign c53ibus[temp_w*4 +:temp_w] = v1212obus[temp_w*0 +:temp_w];
assign v1212ibus[data_w*0 +:data_w] = c53obus[data_w*4 +:data_w];
assign c53ibus[temp_w*5 +:temp_w] = v1301obus[temp_w*0 +:temp_w];
assign v1301ibus[data_w*0 +:data_w] = c53obus[data_w*5 +:data_w];
assign c54ibus[temp_w*0 +:temp_w] = v148obus[temp_w*0 +:temp_w];
assign v148ibus[data_w*0 +:data_w] = c54obus[data_w*0 +:data_w];
assign c54ibus[temp_w*1 +:temp_w] = v223obus[temp_w*0 +:temp_w];
assign v223ibus[data_w*0 +:data_w] = c54obus[data_w*1 +:data_w];
assign c54ibus[temp_w*2 +:temp_w] = v781obus[temp_w*0 +:temp_w];
assign v781ibus[data_w*0 +:data_w] = c54obus[data_w*2 +:data_w];
assign c54ibus[temp_w*3 +:temp_w] = v905obus[temp_w*0 +:temp_w];
assign v905ibus[data_w*0 +:data_w] = c54obus[data_w*3 +:data_w];
assign c54ibus[temp_w*4 +:temp_w] = v1213obus[temp_w*0 +:temp_w];
assign v1213ibus[data_w*0 +:data_w] = c54obus[data_w*4 +:data_w];
assign c54ibus[temp_w*5 +:temp_w] = v1302obus[temp_w*0 +:temp_w];
assign v1302ibus[data_w*0 +:data_w] = c54obus[data_w*5 +:data_w];
assign c55ibus[temp_w*0 +:temp_w] = v149obus[temp_w*0 +:temp_w];
assign v149ibus[data_w*0 +:data_w] = c55obus[data_w*0 +:data_w];
assign c55ibus[temp_w*1 +:temp_w] = v224obus[temp_w*0 +:temp_w];
assign v224ibus[data_w*0 +:data_w] = c55obus[data_w*1 +:data_w];
assign c55ibus[temp_w*2 +:temp_w] = v782obus[temp_w*0 +:temp_w];
assign v782ibus[data_w*0 +:data_w] = c55obus[data_w*2 +:data_w];
assign c55ibus[temp_w*3 +:temp_w] = v906obus[temp_w*0 +:temp_w];
assign v906ibus[data_w*0 +:data_w] = c55obus[data_w*3 +:data_w];
assign c55ibus[temp_w*4 +:temp_w] = v1214obus[temp_w*0 +:temp_w];
assign v1214ibus[data_w*0 +:data_w] = c55obus[data_w*4 +:data_w];
assign c55ibus[temp_w*5 +:temp_w] = v1303obus[temp_w*0 +:temp_w];
assign v1303ibus[data_w*0 +:data_w] = c55obus[data_w*5 +:data_w];
assign c56ibus[temp_w*0 +:temp_w] = v150obus[temp_w*0 +:temp_w];
assign v150ibus[data_w*0 +:data_w] = c56obus[data_w*0 +:data_w];
assign c56ibus[temp_w*1 +:temp_w] = v225obus[temp_w*0 +:temp_w];
assign v225ibus[data_w*0 +:data_w] = c56obus[data_w*1 +:data_w];
assign c56ibus[temp_w*2 +:temp_w] = v783obus[temp_w*0 +:temp_w];
assign v783ibus[data_w*0 +:data_w] = c56obus[data_w*2 +:data_w];
assign c56ibus[temp_w*3 +:temp_w] = v907obus[temp_w*0 +:temp_w];
assign v907ibus[data_w*0 +:data_w] = c56obus[data_w*3 +:data_w];
assign c56ibus[temp_w*4 +:temp_w] = v1215obus[temp_w*0 +:temp_w];
assign v1215ibus[data_w*0 +:data_w] = c56obus[data_w*4 +:data_w];
assign c56ibus[temp_w*5 +:temp_w] = v1304obus[temp_w*0 +:temp_w];
assign v1304ibus[data_w*0 +:data_w] = c56obus[data_w*5 +:data_w];
assign c57ibus[temp_w*0 +:temp_w] = v151obus[temp_w*0 +:temp_w];
assign v151ibus[data_w*0 +:data_w] = c57obus[data_w*0 +:data_w];
assign c57ibus[temp_w*1 +:temp_w] = v226obus[temp_w*0 +:temp_w];
assign v226ibus[data_w*0 +:data_w] = c57obus[data_w*1 +:data_w];
assign c57ibus[temp_w*2 +:temp_w] = v784obus[temp_w*0 +:temp_w];
assign v784ibus[data_w*0 +:data_w] = c57obus[data_w*2 +:data_w];
assign c57ibus[temp_w*3 +:temp_w] = v908obus[temp_w*0 +:temp_w];
assign v908ibus[data_w*0 +:data_w] = c57obus[data_w*3 +:data_w];
assign c57ibus[temp_w*4 +:temp_w] = v1216obus[temp_w*0 +:temp_w];
assign v1216ibus[data_w*0 +:data_w] = c57obus[data_w*4 +:data_w];
assign c57ibus[temp_w*5 +:temp_w] = v1305obus[temp_w*0 +:temp_w];
assign v1305ibus[data_w*0 +:data_w] = c57obus[data_w*5 +:data_w];
assign c58ibus[temp_w*0 +:temp_w] = v152obus[temp_w*0 +:temp_w];
assign v152ibus[data_w*0 +:data_w] = c58obus[data_w*0 +:data_w];
assign c58ibus[temp_w*1 +:temp_w] = v227obus[temp_w*0 +:temp_w];
assign v227ibus[data_w*0 +:data_w] = c58obus[data_w*1 +:data_w];
assign c58ibus[temp_w*2 +:temp_w] = v785obus[temp_w*0 +:temp_w];
assign v785ibus[data_w*0 +:data_w] = c58obus[data_w*2 +:data_w];
assign c58ibus[temp_w*3 +:temp_w] = v909obus[temp_w*0 +:temp_w];
assign v909ibus[data_w*0 +:data_w] = c58obus[data_w*3 +:data_w];
assign c58ibus[temp_w*4 +:temp_w] = v1217obus[temp_w*0 +:temp_w];
assign v1217ibus[data_w*0 +:data_w] = c58obus[data_w*4 +:data_w];
assign c58ibus[temp_w*5 +:temp_w] = v1306obus[temp_w*0 +:temp_w];
assign v1306ibus[data_w*0 +:data_w] = c58obus[data_w*5 +:data_w];
assign c59ibus[temp_w*0 +:temp_w] = v153obus[temp_w*0 +:temp_w];
assign v153ibus[data_w*0 +:data_w] = c59obus[data_w*0 +:data_w];
assign c59ibus[temp_w*1 +:temp_w] = v228obus[temp_w*0 +:temp_w];
assign v228ibus[data_w*0 +:data_w] = c59obus[data_w*1 +:data_w];
assign c59ibus[temp_w*2 +:temp_w] = v786obus[temp_w*0 +:temp_w];
assign v786ibus[data_w*0 +:data_w] = c59obus[data_w*2 +:data_w];
assign c59ibus[temp_w*3 +:temp_w] = v910obus[temp_w*0 +:temp_w];
assign v910ibus[data_w*0 +:data_w] = c59obus[data_w*3 +:data_w];
assign c59ibus[temp_w*4 +:temp_w] = v1218obus[temp_w*0 +:temp_w];
assign v1218ibus[data_w*0 +:data_w] = c59obus[data_w*4 +:data_w];
assign c59ibus[temp_w*5 +:temp_w] = v1307obus[temp_w*0 +:temp_w];
assign v1307ibus[data_w*0 +:data_w] = c59obus[data_w*5 +:data_w];
assign c60ibus[temp_w*0 +:temp_w] = v154obus[temp_w*0 +:temp_w];
assign v154ibus[data_w*0 +:data_w] = c60obus[data_w*0 +:data_w];
assign c60ibus[temp_w*1 +:temp_w] = v229obus[temp_w*0 +:temp_w];
assign v229ibus[data_w*0 +:data_w] = c60obus[data_w*1 +:data_w];
assign c60ibus[temp_w*2 +:temp_w] = v787obus[temp_w*0 +:temp_w];
assign v787ibus[data_w*0 +:data_w] = c60obus[data_w*2 +:data_w];
assign c60ibus[temp_w*3 +:temp_w] = v911obus[temp_w*0 +:temp_w];
assign v911ibus[data_w*0 +:data_w] = c60obus[data_w*3 +:data_w];
assign c60ibus[temp_w*4 +:temp_w] = v1219obus[temp_w*0 +:temp_w];
assign v1219ibus[data_w*0 +:data_w] = c60obus[data_w*4 +:data_w];
assign c60ibus[temp_w*5 +:temp_w] = v1308obus[temp_w*0 +:temp_w];
assign v1308ibus[data_w*0 +:data_w] = c60obus[data_w*5 +:data_w];
assign c61ibus[temp_w*0 +:temp_w] = v155obus[temp_w*0 +:temp_w];
assign v155ibus[data_w*0 +:data_w] = c61obus[data_w*0 +:data_w];
assign c61ibus[temp_w*1 +:temp_w] = v230obus[temp_w*0 +:temp_w];
assign v230ibus[data_w*0 +:data_w] = c61obus[data_w*1 +:data_w];
assign c61ibus[temp_w*2 +:temp_w] = v788obus[temp_w*0 +:temp_w];
assign v788ibus[data_w*0 +:data_w] = c61obus[data_w*2 +:data_w];
assign c61ibus[temp_w*3 +:temp_w] = v912obus[temp_w*0 +:temp_w];
assign v912ibus[data_w*0 +:data_w] = c61obus[data_w*3 +:data_w];
assign c61ibus[temp_w*4 +:temp_w] = v1220obus[temp_w*0 +:temp_w];
assign v1220ibus[data_w*0 +:data_w] = c61obus[data_w*4 +:data_w];
assign c61ibus[temp_w*5 +:temp_w] = v1309obus[temp_w*0 +:temp_w];
assign v1309ibus[data_w*0 +:data_w] = c61obus[data_w*5 +:data_w];
assign c62ibus[temp_w*0 +:temp_w] = v156obus[temp_w*0 +:temp_w];
assign v156ibus[data_w*0 +:data_w] = c62obus[data_w*0 +:data_w];
assign c62ibus[temp_w*1 +:temp_w] = v231obus[temp_w*0 +:temp_w];
assign v231ibus[data_w*0 +:data_w] = c62obus[data_w*1 +:data_w];
assign c62ibus[temp_w*2 +:temp_w] = v789obus[temp_w*0 +:temp_w];
assign v789ibus[data_w*0 +:data_w] = c62obus[data_w*2 +:data_w];
assign c62ibus[temp_w*3 +:temp_w] = v913obus[temp_w*0 +:temp_w];
assign v913ibus[data_w*0 +:data_w] = c62obus[data_w*3 +:data_w];
assign c62ibus[temp_w*4 +:temp_w] = v1221obus[temp_w*0 +:temp_w];
assign v1221ibus[data_w*0 +:data_w] = c62obus[data_w*4 +:data_w];
assign c62ibus[temp_w*5 +:temp_w] = v1310obus[temp_w*0 +:temp_w];
assign v1310ibus[data_w*0 +:data_w] = c62obus[data_w*5 +:data_w];
assign c63ibus[temp_w*0 +:temp_w] = v157obus[temp_w*0 +:temp_w];
assign v157ibus[data_w*0 +:data_w] = c63obus[data_w*0 +:data_w];
assign c63ibus[temp_w*1 +:temp_w] = v232obus[temp_w*0 +:temp_w];
assign v232ibus[data_w*0 +:data_w] = c63obus[data_w*1 +:data_w];
assign c63ibus[temp_w*2 +:temp_w] = v790obus[temp_w*0 +:temp_w];
assign v790ibus[data_w*0 +:data_w] = c63obus[data_w*2 +:data_w];
assign c63ibus[temp_w*3 +:temp_w] = v914obus[temp_w*0 +:temp_w];
assign v914ibus[data_w*0 +:data_w] = c63obus[data_w*3 +:data_w];
assign c63ibus[temp_w*4 +:temp_w] = v1222obus[temp_w*0 +:temp_w];
assign v1222ibus[data_w*0 +:data_w] = c63obus[data_w*4 +:data_w];
assign c63ibus[temp_w*5 +:temp_w] = v1311obus[temp_w*0 +:temp_w];
assign v1311ibus[data_w*0 +:data_w] = c63obus[data_w*5 +:data_w];
assign c64ibus[temp_w*0 +:temp_w] = v158obus[temp_w*0 +:temp_w];
assign v158ibus[data_w*0 +:data_w] = c64obus[data_w*0 +:data_w];
assign c64ibus[temp_w*1 +:temp_w] = v233obus[temp_w*0 +:temp_w];
assign v233ibus[data_w*0 +:data_w] = c64obus[data_w*1 +:data_w];
assign c64ibus[temp_w*2 +:temp_w] = v791obus[temp_w*0 +:temp_w];
assign v791ibus[data_w*0 +:data_w] = c64obus[data_w*2 +:data_w];
assign c64ibus[temp_w*3 +:temp_w] = v915obus[temp_w*0 +:temp_w];
assign v915ibus[data_w*0 +:data_w] = c64obus[data_w*3 +:data_w];
assign c64ibus[temp_w*4 +:temp_w] = v1223obus[temp_w*0 +:temp_w];
assign v1223ibus[data_w*0 +:data_w] = c64obus[data_w*4 +:data_w];
assign c64ibus[temp_w*5 +:temp_w] = v1312obus[temp_w*0 +:temp_w];
assign v1312ibus[data_w*0 +:data_w] = c64obus[data_w*5 +:data_w];
assign c65ibus[temp_w*0 +:temp_w] = v159obus[temp_w*0 +:temp_w];
assign v159ibus[data_w*0 +:data_w] = c65obus[data_w*0 +:data_w];
assign c65ibus[temp_w*1 +:temp_w] = v234obus[temp_w*0 +:temp_w];
assign v234ibus[data_w*0 +:data_w] = c65obus[data_w*1 +:data_w];
assign c65ibus[temp_w*2 +:temp_w] = v792obus[temp_w*0 +:temp_w];
assign v792ibus[data_w*0 +:data_w] = c65obus[data_w*2 +:data_w];
assign c65ibus[temp_w*3 +:temp_w] = v916obus[temp_w*0 +:temp_w];
assign v916ibus[data_w*0 +:data_w] = c65obus[data_w*3 +:data_w];
assign c65ibus[temp_w*4 +:temp_w] = v1224obus[temp_w*0 +:temp_w];
assign v1224ibus[data_w*0 +:data_w] = c65obus[data_w*4 +:data_w];
assign c65ibus[temp_w*5 +:temp_w] = v1313obus[temp_w*0 +:temp_w];
assign v1313ibus[data_w*0 +:data_w] = c65obus[data_w*5 +:data_w];
assign c66ibus[temp_w*0 +:temp_w] = v160obus[temp_w*0 +:temp_w];
assign v160ibus[data_w*0 +:data_w] = c66obus[data_w*0 +:data_w];
assign c66ibus[temp_w*1 +:temp_w] = v235obus[temp_w*0 +:temp_w];
assign v235ibus[data_w*0 +:data_w] = c66obus[data_w*1 +:data_w];
assign c66ibus[temp_w*2 +:temp_w] = v793obus[temp_w*0 +:temp_w];
assign v793ibus[data_w*0 +:data_w] = c66obus[data_w*2 +:data_w];
assign c66ibus[temp_w*3 +:temp_w] = v917obus[temp_w*0 +:temp_w];
assign v917ibus[data_w*0 +:data_w] = c66obus[data_w*3 +:data_w];
assign c66ibus[temp_w*4 +:temp_w] = v1225obus[temp_w*0 +:temp_w];
assign v1225ibus[data_w*0 +:data_w] = c66obus[data_w*4 +:data_w];
assign c66ibus[temp_w*5 +:temp_w] = v1314obus[temp_w*0 +:temp_w];
assign v1314ibus[data_w*0 +:data_w] = c66obus[data_w*5 +:data_w];
assign c67ibus[temp_w*0 +:temp_w] = v161obus[temp_w*0 +:temp_w];
assign v161ibus[data_w*0 +:data_w] = c67obus[data_w*0 +:data_w];
assign c67ibus[temp_w*1 +:temp_w] = v236obus[temp_w*0 +:temp_w];
assign v236ibus[data_w*0 +:data_w] = c67obus[data_w*1 +:data_w];
assign c67ibus[temp_w*2 +:temp_w] = v794obus[temp_w*0 +:temp_w];
assign v794ibus[data_w*0 +:data_w] = c67obus[data_w*2 +:data_w];
assign c67ibus[temp_w*3 +:temp_w] = v918obus[temp_w*0 +:temp_w];
assign v918ibus[data_w*0 +:data_w] = c67obus[data_w*3 +:data_w];
assign c67ibus[temp_w*4 +:temp_w] = v1226obus[temp_w*0 +:temp_w];
assign v1226ibus[data_w*0 +:data_w] = c67obus[data_w*4 +:data_w];
assign c67ibus[temp_w*5 +:temp_w] = v1315obus[temp_w*0 +:temp_w];
assign v1315ibus[data_w*0 +:data_w] = c67obus[data_w*5 +:data_w];
assign c68ibus[temp_w*0 +:temp_w] = v162obus[temp_w*0 +:temp_w];
assign v162ibus[data_w*0 +:data_w] = c68obus[data_w*0 +:data_w];
assign c68ibus[temp_w*1 +:temp_w] = v237obus[temp_w*0 +:temp_w];
assign v237ibus[data_w*0 +:data_w] = c68obus[data_w*1 +:data_w];
assign c68ibus[temp_w*2 +:temp_w] = v795obus[temp_w*0 +:temp_w];
assign v795ibus[data_w*0 +:data_w] = c68obus[data_w*2 +:data_w];
assign c68ibus[temp_w*3 +:temp_w] = v919obus[temp_w*0 +:temp_w];
assign v919ibus[data_w*0 +:data_w] = c68obus[data_w*3 +:data_w];
assign c68ibus[temp_w*4 +:temp_w] = v1227obus[temp_w*0 +:temp_w];
assign v1227ibus[data_w*0 +:data_w] = c68obus[data_w*4 +:data_w];
assign c68ibus[temp_w*5 +:temp_w] = v1316obus[temp_w*0 +:temp_w];
assign v1316ibus[data_w*0 +:data_w] = c68obus[data_w*5 +:data_w];
assign c69ibus[temp_w*0 +:temp_w] = v163obus[temp_w*0 +:temp_w];
assign v163ibus[data_w*0 +:data_w] = c69obus[data_w*0 +:data_w];
assign c69ibus[temp_w*1 +:temp_w] = v238obus[temp_w*0 +:temp_w];
assign v238ibus[data_w*0 +:data_w] = c69obus[data_w*1 +:data_w];
assign c69ibus[temp_w*2 +:temp_w] = v796obus[temp_w*0 +:temp_w];
assign v796ibus[data_w*0 +:data_w] = c69obus[data_w*2 +:data_w];
assign c69ibus[temp_w*3 +:temp_w] = v920obus[temp_w*0 +:temp_w];
assign v920ibus[data_w*0 +:data_w] = c69obus[data_w*3 +:data_w];
assign c69ibus[temp_w*4 +:temp_w] = v1228obus[temp_w*0 +:temp_w];
assign v1228ibus[data_w*0 +:data_w] = c69obus[data_w*4 +:data_w];
assign c69ibus[temp_w*5 +:temp_w] = v1317obus[temp_w*0 +:temp_w];
assign v1317ibus[data_w*0 +:data_w] = c69obus[data_w*5 +:data_w];
assign c70ibus[temp_w*0 +:temp_w] = v164obus[temp_w*0 +:temp_w];
assign v164ibus[data_w*0 +:data_w] = c70obus[data_w*0 +:data_w];
assign c70ibus[temp_w*1 +:temp_w] = v239obus[temp_w*0 +:temp_w];
assign v239ibus[data_w*0 +:data_w] = c70obus[data_w*1 +:data_w];
assign c70ibus[temp_w*2 +:temp_w] = v797obus[temp_w*0 +:temp_w];
assign v797ibus[data_w*0 +:data_w] = c70obus[data_w*2 +:data_w];
assign c70ibus[temp_w*3 +:temp_w] = v921obus[temp_w*0 +:temp_w];
assign v921ibus[data_w*0 +:data_w] = c70obus[data_w*3 +:data_w];
assign c70ibus[temp_w*4 +:temp_w] = v1229obus[temp_w*0 +:temp_w];
assign v1229ibus[data_w*0 +:data_w] = c70obus[data_w*4 +:data_w];
assign c70ibus[temp_w*5 +:temp_w] = v1318obus[temp_w*0 +:temp_w];
assign v1318ibus[data_w*0 +:data_w] = c70obus[data_w*5 +:data_w];
assign c71ibus[temp_w*0 +:temp_w] = v165obus[temp_w*0 +:temp_w];
assign v165ibus[data_w*0 +:data_w] = c71obus[data_w*0 +:data_w];
assign c71ibus[temp_w*1 +:temp_w] = v240obus[temp_w*0 +:temp_w];
assign v240ibus[data_w*0 +:data_w] = c71obus[data_w*1 +:data_w];
assign c71ibus[temp_w*2 +:temp_w] = v798obus[temp_w*0 +:temp_w];
assign v798ibus[data_w*0 +:data_w] = c71obus[data_w*2 +:data_w];
assign c71ibus[temp_w*3 +:temp_w] = v922obus[temp_w*0 +:temp_w];
assign v922ibus[data_w*0 +:data_w] = c71obus[data_w*3 +:data_w];
assign c71ibus[temp_w*4 +:temp_w] = v1230obus[temp_w*0 +:temp_w];
assign v1230ibus[data_w*0 +:data_w] = c71obus[data_w*4 +:data_w];
assign c71ibus[temp_w*5 +:temp_w] = v1319obus[temp_w*0 +:temp_w];
assign v1319ibus[data_w*0 +:data_w] = c71obus[data_w*5 +:data_w];
assign c72ibus[temp_w*0 +:temp_w] = v166obus[temp_w*0 +:temp_w];
assign v166ibus[data_w*0 +:data_w] = c72obus[data_w*0 +:data_w];
assign c72ibus[temp_w*1 +:temp_w] = v241obus[temp_w*0 +:temp_w];
assign v241ibus[data_w*0 +:data_w] = c72obus[data_w*1 +:data_w];
assign c72ibus[temp_w*2 +:temp_w] = v799obus[temp_w*0 +:temp_w];
assign v799ibus[data_w*0 +:data_w] = c72obus[data_w*2 +:data_w];
assign c72ibus[temp_w*3 +:temp_w] = v923obus[temp_w*0 +:temp_w];
assign v923ibus[data_w*0 +:data_w] = c72obus[data_w*3 +:data_w];
assign c72ibus[temp_w*4 +:temp_w] = v1231obus[temp_w*0 +:temp_w];
assign v1231ibus[data_w*0 +:data_w] = c72obus[data_w*4 +:data_w];
assign c72ibus[temp_w*5 +:temp_w] = v1320obus[temp_w*0 +:temp_w];
assign v1320ibus[data_w*0 +:data_w] = c72obus[data_w*5 +:data_w];
assign c73ibus[temp_w*0 +:temp_w] = v167obus[temp_w*0 +:temp_w];
assign v167ibus[data_w*0 +:data_w] = c73obus[data_w*0 +:data_w];
assign c73ibus[temp_w*1 +:temp_w] = v242obus[temp_w*0 +:temp_w];
assign v242ibus[data_w*0 +:data_w] = c73obus[data_w*1 +:data_w];
assign c73ibus[temp_w*2 +:temp_w] = v800obus[temp_w*0 +:temp_w];
assign v800ibus[data_w*0 +:data_w] = c73obus[data_w*2 +:data_w];
assign c73ibus[temp_w*3 +:temp_w] = v924obus[temp_w*0 +:temp_w];
assign v924ibus[data_w*0 +:data_w] = c73obus[data_w*3 +:data_w];
assign c73ibus[temp_w*4 +:temp_w] = v1232obus[temp_w*0 +:temp_w];
assign v1232ibus[data_w*0 +:data_w] = c73obus[data_w*4 +:data_w];
assign c73ibus[temp_w*5 +:temp_w] = v1321obus[temp_w*0 +:temp_w];
assign v1321ibus[data_w*0 +:data_w] = c73obus[data_w*5 +:data_w];
assign c74ibus[temp_w*0 +:temp_w] = v168obus[temp_w*0 +:temp_w];
assign v168ibus[data_w*0 +:data_w] = c74obus[data_w*0 +:data_w];
assign c74ibus[temp_w*1 +:temp_w] = v243obus[temp_w*0 +:temp_w];
assign v243ibus[data_w*0 +:data_w] = c74obus[data_w*1 +:data_w];
assign c74ibus[temp_w*2 +:temp_w] = v801obus[temp_w*0 +:temp_w];
assign v801ibus[data_w*0 +:data_w] = c74obus[data_w*2 +:data_w];
assign c74ibus[temp_w*3 +:temp_w] = v925obus[temp_w*0 +:temp_w];
assign v925ibus[data_w*0 +:data_w] = c74obus[data_w*3 +:data_w];
assign c74ibus[temp_w*4 +:temp_w] = v1233obus[temp_w*0 +:temp_w];
assign v1233ibus[data_w*0 +:data_w] = c74obus[data_w*4 +:data_w];
assign c74ibus[temp_w*5 +:temp_w] = v1322obus[temp_w*0 +:temp_w];
assign v1322ibus[data_w*0 +:data_w] = c74obus[data_w*5 +:data_w];
assign c75ibus[temp_w*0 +:temp_w] = v169obus[temp_w*0 +:temp_w];
assign v169ibus[data_w*0 +:data_w] = c75obus[data_w*0 +:data_w];
assign c75ibus[temp_w*1 +:temp_w] = v244obus[temp_w*0 +:temp_w];
assign v244ibus[data_w*0 +:data_w] = c75obus[data_w*1 +:data_w];
assign c75ibus[temp_w*2 +:temp_w] = v802obus[temp_w*0 +:temp_w];
assign v802ibus[data_w*0 +:data_w] = c75obus[data_w*2 +:data_w];
assign c75ibus[temp_w*3 +:temp_w] = v926obus[temp_w*0 +:temp_w];
assign v926ibus[data_w*0 +:data_w] = c75obus[data_w*3 +:data_w];
assign c75ibus[temp_w*4 +:temp_w] = v1234obus[temp_w*0 +:temp_w];
assign v1234ibus[data_w*0 +:data_w] = c75obus[data_w*4 +:data_w];
assign c75ibus[temp_w*5 +:temp_w] = v1323obus[temp_w*0 +:temp_w];
assign v1323ibus[data_w*0 +:data_w] = c75obus[data_w*5 +:data_w];
assign c76ibus[temp_w*0 +:temp_w] = v170obus[temp_w*0 +:temp_w];
assign v170ibus[data_w*0 +:data_w] = c76obus[data_w*0 +:data_w];
assign c76ibus[temp_w*1 +:temp_w] = v245obus[temp_w*0 +:temp_w];
assign v245ibus[data_w*0 +:data_w] = c76obus[data_w*1 +:data_w];
assign c76ibus[temp_w*2 +:temp_w] = v803obus[temp_w*0 +:temp_w];
assign v803ibus[data_w*0 +:data_w] = c76obus[data_w*2 +:data_w];
assign c76ibus[temp_w*3 +:temp_w] = v927obus[temp_w*0 +:temp_w];
assign v927ibus[data_w*0 +:data_w] = c76obus[data_w*3 +:data_w];
assign c76ibus[temp_w*4 +:temp_w] = v1235obus[temp_w*0 +:temp_w];
assign v1235ibus[data_w*0 +:data_w] = c76obus[data_w*4 +:data_w];
assign c76ibus[temp_w*5 +:temp_w] = v1324obus[temp_w*0 +:temp_w];
assign v1324ibus[data_w*0 +:data_w] = c76obus[data_w*5 +:data_w];
assign c77ibus[temp_w*0 +:temp_w] = v171obus[temp_w*0 +:temp_w];
assign v171ibus[data_w*0 +:data_w] = c77obus[data_w*0 +:data_w];
assign c77ibus[temp_w*1 +:temp_w] = v246obus[temp_w*0 +:temp_w];
assign v246ibus[data_w*0 +:data_w] = c77obus[data_w*1 +:data_w];
assign c77ibus[temp_w*2 +:temp_w] = v804obus[temp_w*0 +:temp_w];
assign v804ibus[data_w*0 +:data_w] = c77obus[data_w*2 +:data_w];
assign c77ibus[temp_w*3 +:temp_w] = v928obus[temp_w*0 +:temp_w];
assign v928ibus[data_w*0 +:data_w] = c77obus[data_w*3 +:data_w];
assign c77ibus[temp_w*4 +:temp_w] = v1236obus[temp_w*0 +:temp_w];
assign v1236ibus[data_w*0 +:data_w] = c77obus[data_w*4 +:data_w];
assign c77ibus[temp_w*5 +:temp_w] = v1325obus[temp_w*0 +:temp_w];
assign v1325ibus[data_w*0 +:data_w] = c77obus[data_w*5 +:data_w];
assign c78ibus[temp_w*0 +:temp_w] = v172obus[temp_w*0 +:temp_w];
assign v172ibus[data_w*0 +:data_w] = c78obus[data_w*0 +:data_w];
assign c78ibus[temp_w*1 +:temp_w] = v247obus[temp_w*0 +:temp_w];
assign v247ibus[data_w*0 +:data_w] = c78obus[data_w*1 +:data_w];
assign c78ibus[temp_w*2 +:temp_w] = v805obus[temp_w*0 +:temp_w];
assign v805ibus[data_w*0 +:data_w] = c78obus[data_w*2 +:data_w];
assign c78ibus[temp_w*3 +:temp_w] = v929obus[temp_w*0 +:temp_w];
assign v929ibus[data_w*0 +:data_w] = c78obus[data_w*3 +:data_w];
assign c78ibus[temp_w*4 +:temp_w] = v1237obus[temp_w*0 +:temp_w];
assign v1237ibus[data_w*0 +:data_w] = c78obus[data_w*4 +:data_w];
assign c78ibus[temp_w*5 +:temp_w] = v1326obus[temp_w*0 +:temp_w];
assign v1326ibus[data_w*0 +:data_w] = c78obus[data_w*5 +:data_w];
assign c79ibus[temp_w*0 +:temp_w] = v173obus[temp_w*0 +:temp_w];
assign v173ibus[data_w*0 +:data_w] = c79obus[data_w*0 +:data_w];
assign c79ibus[temp_w*1 +:temp_w] = v248obus[temp_w*0 +:temp_w];
assign v248ibus[data_w*0 +:data_w] = c79obus[data_w*1 +:data_w];
assign c79ibus[temp_w*2 +:temp_w] = v806obus[temp_w*0 +:temp_w];
assign v806ibus[data_w*0 +:data_w] = c79obus[data_w*2 +:data_w];
assign c79ibus[temp_w*3 +:temp_w] = v930obus[temp_w*0 +:temp_w];
assign v930ibus[data_w*0 +:data_w] = c79obus[data_w*3 +:data_w];
assign c79ibus[temp_w*4 +:temp_w] = v1238obus[temp_w*0 +:temp_w];
assign v1238ibus[data_w*0 +:data_w] = c79obus[data_w*4 +:data_w];
assign c79ibus[temp_w*5 +:temp_w] = v1327obus[temp_w*0 +:temp_w];
assign v1327ibus[data_w*0 +:data_w] = c79obus[data_w*5 +:data_w];
assign c80ibus[temp_w*0 +:temp_w] = v174obus[temp_w*0 +:temp_w];
assign v174ibus[data_w*0 +:data_w] = c80obus[data_w*0 +:data_w];
assign c80ibus[temp_w*1 +:temp_w] = v249obus[temp_w*0 +:temp_w];
assign v249ibus[data_w*0 +:data_w] = c80obus[data_w*1 +:data_w];
assign c80ibus[temp_w*2 +:temp_w] = v807obus[temp_w*0 +:temp_w];
assign v807ibus[data_w*0 +:data_w] = c80obus[data_w*2 +:data_w];
assign c80ibus[temp_w*3 +:temp_w] = v931obus[temp_w*0 +:temp_w];
assign v931ibus[data_w*0 +:data_w] = c80obus[data_w*3 +:data_w];
assign c80ibus[temp_w*4 +:temp_w] = v1239obus[temp_w*0 +:temp_w];
assign v1239ibus[data_w*0 +:data_w] = c80obus[data_w*4 +:data_w];
assign c80ibus[temp_w*5 +:temp_w] = v1328obus[temp_w*0 +:temp_w];
assign v1328ibus[data_w*0 +:data_w] = c80obus[data_w*5 +:data_w];
assign c81ibus[temp_w*0 +:temp_w] = v175obus[temp_w*0 +:temp_w];
assign v175ibus[data_w*0 +:data_w] = c81obus[data_w*0 +:data_w];
assign c81ibus[temp_w*1 +:temp_w] = v250obus[temp_w*0 +:temp_w];
assign v250ibus[data_w*0 +:data_w] = c81obus[data_w*1 +:data_w];
assign c81ibus[temp_w*2 +:temp_w] = v808obus[temp_w*0 +:temp_w];
assign v808ibus[data_w*0 +:data_w] = c81obus[data_w*2 +:data_w];
assign c81ibus[temp_w*3 +:temp_w] = v932obus[temp_w*0 +:temp_w];
assign v932ibus[data_w*0 +:data_w] = c81obus[data_w*3 +:data_w];
assign c81ibus[temp_w*4 +:temp_w] = v1240obus[temp_w*0 +:temp_w];
assign v1240ibus[data_w*0 +:data_w] = c81obus[data_w*4 +:data_w];
assign c81ibus[temp_w*5 +:temp_w] = v1329obus[temp_w*0 +:temp_w];
assign v1329ibus[data_w*0 +:data_w] = c81obus[data_w*5 +:data_w];
assign c82ibus[temp_w*0 +:temp_w] = v176obus[temp_w*0 +:temp_w];
assign v176ibus[data_w*0 +:data_w] = c82obus[data_w*0 +:data_w];
assign c82ibus[temp_w*1 +:temp_w] = v251obus[temp_w*0 +:temp_w];
assign v251ibus[data_w*0 +:data_w] = c82obus[data_w*1 +:data_w];
assign c82ibus[temp_w*2 +:temp_w] = v809obus[temp_w*0 +:temp_w];
assign v809ibus[data_w*0 +:data_w] = c82obus[data_w*2 +:data_w];
assign c82ibus[temp_w*3 +:temp_w] = v933obus[temp_w*0 +:temp_w];
assign v933ibus[data_w*0 +:data_w] = c82obus[data_w*3 +:data_w];
assign c82ibus[temp_w*4 +:temp_w] = v1241obus[temp_w*0 +:temp_w];
assign v1241ibus[data_w*0 +:data_w] = c82obus[data_w*4 +:data_w];
assign c82ibus[temp_w*5 +:temp_w] = v1330obus[temp_w*0 +:temp_w];
assign v1330ibus[data_w*0 +:data_w] = c82obus[data_w*5 +:data_w];
assign c83ibus[temp_w*0 +:temp_w] = v177obus[temp_w*0 +:temp_w];
assign v177ibus[data_w*0 +:data_w] = c83obus[data_w*0 +:data_w];
assign c83ibus[temp_w*1 +:temp_w] = v252obus[temp_w*0 +:temp_w];
assign v252ibus[data_w*0 +:data_w] = c83obus[data_w*1 +:data_w];
assign c83ibus[temp_w*2 +:temp_w] = v810obus[temp_w*0 +:temp_w];
assign v810ibus[data_w*0 +:data_w] = c83obus[data_w*2 +:data_w];
assign c83ibus[temp_w*3 +:temp_w] = v934obus[temp_w*0 +:temp_w];
assign v934ibus[data_w*0 +:data_w] = c83obus[data_w*3 +:data_w];
assign c83ibus[temp_w*4 +:temp_w] = v1242obus[temp_w*0 +:temp_w];
assign v1242ibus[data_w*0 +:data_w] = c83obus[data_w*4 +:data_w];
assign c83ibus[temp_w*5 +:temp_w] = v1331obus[temp_w*0 +:temp_w];
assign v1331ibus[data_w*0 +:data_w] = c83obus[data_w*5 +:data_w];
assign c84ibus[temp_w*0 +:temp_w] = v178obus[temp_w*0 +:temp_w];
assign v178ibus[data_w*0 +:data_w] = c84obus[data_w*0 +:data_w];
assign c84ibus[temp_w*1 +:temp_w] = v253obus[temp_w*0 +:temp_w];
assign v253ibus[data_w*0 +:data_w] = c84obus[data_w*1 +:data_w];
assign c84ibus[temp_w*2 +:temp_w] = v811obus[temp_w*0 +:temp_w];
assign v811ibus[data_w*0 +:data_w] = c84obus[data_w*2 +:data_w];
assign c84ibus[temp_w*3 +:temp_w] = v935obus[temp_w*0 +:temp_w];
assign v935ibus[data_w*0 +:data_w] = c84obus[data_w*3 +:data_w];
assign c84ibus[temp_w*4 +:temp_w] = v1243obus[temp_w*0 +:temp_w];
assign v1243ibus[data_w*0 +:data_w] = c84obus[data_w*4 +:data_w];
assign c84ibus[temp_w*5 +:temp_w] = v1332obus[temp_w*0 +:temp_w];
assign v1332ibus[data_w*0 +:data_w] = c84obus[data_w*5 +:data_w];
assign c85ibus[temp_w*0 +:temp_w] = v179obus[temp_w*0 +:temp_w];
assign v179ibus[data_w*0 +:data_w] = c85obus[data_w*0 +:data_w];
assign c85ibus[temp_w*1 +:temp_w] = v254obus[temp_w*0 +:temp_w];
assign v254ibus[data_w*0 +:data_w] = c85obus[data_w*1 +:data_w];
assign c85ibus[temp_w*2 +:temp_w] = v812obus[temp_w*0 +:temp_w];
assign v812ibus[data_w*0 +:data_w] = c85obus[data_w*2 +:data_w];
assign c85ibus[temp_w*3 +:temp_w] = v936obus[temp_w*0 +:temp_w];
assign v936ibus[data_w*0 +:data_w] = c85obus[data_w*3 +:data_w];
assign c85ibus[temp_w*4 +:temp_w] = v1244obus[temp_w*0 +:temp_w];
assign v1244ibus[data_w*0 +:data_w] = c85obus[data_w*4 +:data_w];
assign c85ibus[temp_w*5 +:temp_w] = v1333obus[temp_w*0 +:temp_w];
assign v1333ibus[data_w*0 +:data_w] = c85obus[data_w*5 +:data_w];
assign c86ibus[temp_w*0 +:temp_w] = v180obus[temp_w*0 +:temp_w];
assign v180ibus[data_w*0 +:data_w] = c86obus[data_w*0 +:data_w];
assign c86ibus[temp_w*1 +:temp_w] = v255obus[temp_w*0 +:temp_w];
assign v255ibus[data_w*0 +:data_w] = c86obus[data_w*1 +:data_w];
assign c86ibus[temp_w*2 +:temp_w] = v813obus[temp_w*0 +:temp_w];
assign v813ibus[data_w*0 +:data_w] = c86obus[data_w*2 +:data_w];
assign c86ibus[temp_w*3 +:temp_w] = v937obus[temp_w*0 +:temp_w];
assign v937ibus[data_w*0 +:data_w] = c86obus[data_w*3 +:data_w];
assign c86ibus[temp_w*4 +:temp_w] = v1245obus[temp_w*0 +:temp_w];
assign v1245ibus[data_w*0 +:data_w] = c86obus[data_w*4 +:data_w];
assign c86ibus[temp_w*5 +:temp_w] = v1334obus[temp_w*0 +:temp_w];
assign v1334ibus[data_w*0 +:data_w] = c86obus[data_w*5 +:data_w];
assign c87ibus[temp_w*0 +:temp_w] = v181obus[temp_w*0 +:temp_w];
assign v181ibus[data_w*0 +:data_w] = c87obus[data_w*0 +:data_w];
assign c87ibus[temp_w*1 +:temp_w] = v256obus[temp_w*0 +:temp_w];
assign v256ibus[data_w*0 +:data_w] = c87obus[data_w*1 +:data_w];
assign c87ibus[temp_w*2 +:temp_w] = v814obus[temp_w*0 +:temp_w];
assign v814ibus[data_w*0 +:data_w] = c87obus[data_w*2 +:data_w];
assign c87ibus[temp_w*3 +:temp_w] = v938obus[temp_w*0 +:temp_w];
assign v938ibus[data_w*0 +:data_w] = c87obus[data_w*3 +:data_w];
assign c87ibus[temp_w*4 +:temp_w] = v1246obus[temp_w*0 +:temp_w];
assign v1246ibus[data_w*0 +:data_w] = c87obus[data_w*4 +:data_w];
assign c87ibus[temp_w*5 +:temp_w] = v1335obus[temp_w*0 +:temp_w];
assign v1335ibus[data_w*0 +:data_w] = c87obus[data_w*5 +:data_w];
assign c88ibus[temp_w*0 +:temp_w] = v182obus[temp_w*0 +:temp_w];
assign v182ibus[data_w*0 +:data_w] = c88obus[data_w*0 +:data_w];
assign c88ibus[temp_w*1 +:temp_w] = v257obus[temp_w*0 +:temp_w];
assign v257ibus[data_w*0 +:data_w] = c88obus[data_w*1 +:data_w];
assign c88ibus[temp_w*2 +:temp_w] = v815obus[temp_w*0 +:temp_w];
assign v815ibus[data_w*0 +:data_w] = c88obus[data_w*2 +:data_w];
assign c88ibus[temp_w*3 +:temp_w] = v939obus[temp_w*0 +:temp_w];
assign v939ibus[data_w*0 +:data_w] = c88obus[data_w*3 +:data_w];
assign c88ibus[temp_w*4 +:temp_w] = v1247obus[temp_w*0 +:temp_w];
assign v1247ibus[data_w*0 +:data_w] = c88obus[data_w*4 +:data_w];
assign c88ibus[temp_w*5 +:temp_w] = v1336obus[temp_w*0 +:temp_w];
assign v1336ibus[data_w*0 +:data_w] = c88obus[data_w*5 +:data_w];
assign c89ibus[temp_w*0 +:temp_w] = v183obus[temp_w*0 +:temp_w];
assign v183ibus[data_w*0 +:data_w] = c89obus[data_w*0 +:data_w];
assign c89ibus[temp_w*1 +:temp_w] = v258obus[temp_w*0 +:temp_w];
assign v258ibus[data_w*0 +:data_w] = c89obus[data_w*1 +:data_w];
assign c89ibus[temp_w*2 +:temp_w] = v816obus[temp_w*0 +:temp_w];
assign v816ibus[data_w*0 +:data_w] = c89obus[data_w*2 +:data_w];
assign c89ibus[temp_w*3 +:temp_w] = v940obus[temp_w*0 +:temp_w];
assign v940ibus[data_w*0 +:data_w] = c89obus[data_w*3 +:data_w];
assign c89ibus[temp_w*4 +:temp_w] = v1152obus[temp_w*0 +:temp_w];
assign v1152ibus[data_w*0 +:data_w] = c89obus[data_w*4 +:data_w];
assign c89ibus[temp_w*5 +:temp_w] = v1337obus[temp_w*0 +:temp_w];
assign v1337ibus[data_w*0 +:data_w] = c89obus[data_w*5 +:data_w];
assign c90ibus[temp_w*0 +:temp_w] = v184obus[temp_w*0 +:temp_w];
assign v184ibus[data_w*0 +:data_w] = c90obus[data_w*0 +:data_w];
assign c90ibus[temp_w*1 +:temp_w] = v259obus[temp_w*0 +:temp_w];
assign v259ibus[data_w*0 +:data_w] = c90obus[data_w*1 +:data_w];
assign c90ibus[temp_w*2 +:temp_w] = v817obus[temp_w*0 +:temp_w];
assign v817ibus[data_w*0 +:data_w] = c90obus[data_w*2 +:data_w];
assign c90ibus[temp_w*3 +:temp_w] = v941obus[temp_w*0 +:temp_w];
assign v941ibus[data_w*0 +:data_w] = c90obus[data_w*3 +:data_w];
assign c90ibus[temp_w*4 +:temp_w] = v1153obus[temp_w*0 +:temp_w];
assign v1153ibus[data_w*0 +:data_w] = c90obus[data_w*4 +:data_w];
assign c90ibus[temp_w*5 +:temp_w] = v1338obus[temp_w*0 +:temp_w];
assign v1338ibus[data_w*0 +:data_w] = c90obus[data_w*5 +:data_w];
assign c91ibus[temp_w*0 +:temp_w] = v185obus[temp_w*0 +:temp_w];
assign v185ibus[data_w*0 +:data_w] = c91obus[data_w*0 +:data_w];
assign c91ibus[temp_w*1 +:temp_w] = v260obus[temp_w*0 +:temp_w];
assign v260ibus[data_w*0 +:data_w] = c91obus[data_w*1 +:data_w];
assign c91ibus[temp_w*2 +:temp_w] = v818obus[temp_w*0 +:temp_w];
assign v818ibus[data_w*0 +:data_w] = c91obus[data_w*2 +:data_w];
assign c91ibus[temp_w*3 +:temp_w] = v942obus[temp_w*0 +:temp_w];
assign v942ibus[data_w*0 +:data_w] = c91obus[data_w*3 +:data_w];
assign c91ibus[temp_w*4 +:temp_w] = v1154obus[temp_w*0 +:temp_w];
assign v1154ibus[data_w*0 +:data_w] = c91obus[data_w*4 +:data_w];
assign c91ibus[temp_w*5 +:temp_w] = v1339obus[temp_w*0 +:temp_w];
assign v1339ibus[data_w*0 +:data_w] = c91obus[data_w*5 +:data_w];
assign c92ibus[temp_w*0 +:temp_w] = v186obus[temp_w*0 +:temp_w];
assign v186ibus[data_w*0 +:data_w] = c92obus[data_w*0 +:data_w];
assign c92ibus[temp_w*1 +:temp_w] = v261obus[temp_w*0 +:temp_w];
assign v261ibus[data_w*0 +:data_w] = c92obus[data_w*1 +:data_w];
assign c92ibus[temp_w*2 +:temp_w] = v819obus[temp_w*0 +:temp_w];
assign v819ibus[data_w*0 +:data_w] = c92obus[data_w*2 +:data_w];
assign c92ibus[temp_w*3 +:temp_w] = v943obus[temp_w*0 +:temp_w];
assign v943ibus[data_w*0 +:data_w] = c92obus[data_w*3 +:data_w];
assign c92ibus[temp_w*4 +:temp_w] = v1155obus[temp_w*0 +:temp_w];
assign v1155ibus[data_w*0 +:data_w] = c92obus[data_w*4 +:data_w];
assign c92ibus[temp_w*5 +:temp_w] = v1340obus[temp_w*0 +:temp_w];
assign v1340ibus[data_w*0 +:data_w] = c92obus[data_w*5 +:data_w];
assign c93ibus[temp_w*0 +:temp_w] = v187obus[temp_w*0 +:temp_w];
assign v187ibus[data_w*0 +:data_w] = c93obus[data_w*0 +:data_w];
assign c93ibus[temp_w*1 +:temp_w] = v262obus[temp_w*0 +:temp_w];
assign v262ibus[data_w*0 +:data_w] = c93obus[data_w*1 +:data_w];
assign c93ibus[temp_w*2 +:temp_w] = v820obus[temp_w*0 +:temp_w];
assign v820ibus[data_w*0 +:data_w] = c93obus[data_w*2 +:data_w];
assign c93ibus[temp_w*3 +:temp_w] = v944obus[temp_w*0 +:temp_w];
assign v944ibus[data_w*0 +:data_w] = c93obus[data_w*3 +:data_w];
assign c93ibus[temp_w*4 +:temp_w] = v1156obus[temp_w*0 +:temp_w];
assign v1156ibus[data_w*0 +:data_w] = c93obus[data_w*4 +:data_w];
assign c93ibus[temp_w*5 +:temp_w] = v1341obus[temp_w*0 +:temp_w];
assign v1341ibus[data_w*0 +:data_w] = c93obus[data_w*5 +:data_w];
assign c94ibus[temp_w*0 +:temp_w] = v188obus[temp_w*0 +:temp_w];
assign v188ibus[data_w*0 +:data_w] = c94obus[data_w*0 +:data_w];
assign c94ibus[temp_w*1 +:temp_w] = v263obus[temp_w*0 +:temp_w];
assign v263ibus[data_w*0 +:data_w] = c94obus[data_w*1 +:data_w];
assign c94ibus[temp_w*2 +:temp_w] = v821obus[temp_w*0 +:temp_w];
assign v821ibus[data_w*0 +:data_w] = c94obus[data_w*2 +:data_w];
assign c94ibus[temp_w*3 +:temp_w] = v945obus[temp_w*0 +:temp_w];
assign v945ibus[data_w*0 +:data_w] = c94obus[data_w*3 +:data_w];
assign c94ibus[temp_w*4 +:temp_w] = v1157obus[temp_w*0 +:temp_w];
assign v1157ibus[data_w*0 +:data_w] = c94obus[data_w*4 +:data_w];
assign c94ibus[temp_w*5 +:temp_w] = v1342obus[temp_w*0 +:temp_w];
assign v1342ibus[data_w*0 +:data_w] = c94obus[data_w*5 +:data_w];
assign c95ibus[temp_w*0 +:temp_w] = v189obus[temp_w*0 +:temp_w];
assign v189ibus[data_w*0 +:data_w] = c95obus[data_w*0 +:data_w];
assign c95ibus[temp_w*1 +:temp_w] = v264obus[temp_w*0 +:temp_w];
assign v264ibus[data_w*0 +:data_w] = c95obus[data_w*1 +:data_w];
assign c95ibus[temp_w*2 +:temp_w] = v822obus[temp_w*0 +:temp_w];
assign v822ibus[data_w*0 +:data_w] = c95obus[data_w*2 +:data_w];
assign c95ibus[temp_w*3 +:temp_w] = v946obus[temp_w*0 +:temp_w];
assign v946ibus[data_w*0 +:data_w] = c95obus[data_w*3 +:data_w];
assign c95ibus[temp_w*4 +:temp_w] = v1158obus[temp_w*0 +:temp_w];
assign v1158ibus[data_w*0 +:data_w] = c95obus[data_w*4 +:data_w];
assign c95ibus[temp_w*5 +:temp_w] = v1343obus[temp_w*0 +:temp_w];
assign v1343ibus[data_w*0 +:data_w] = c95obus[data_w*5 +:data_w];
assign c96ibus[temp_w*0 +:temp_w] = v123obus[temp_w*1 +:temp_w];
assign v123ibus[data_w*1 +:data_w] = c96obus[data_w*0 +:data_w];
assign c96ibus[temp_w*1 +:temp_w] = v502obus[temp_w*0 +:temp_w];
assign v502ibus[data_w*0 +:data_w] = c96obus[data_w*1 +:data_w];
assign c96ibus[temp_w*2 +:temp_w] = v655obus[temp_w*0 +:temp_w];
assign v655ibus[data_w*0 +:data_w] = c96obus[data_w*2 +:data_w];
assign c96ibus[temp_w*3 +:temp_w] = v681obus[temp_w*0 +:temp_w];
assign v681ibus[data_w*0 +:data_w] = c96obus[data_w*3 +:data_w];
assign c96ibus[temp_w*4 +:temp_w] = v1068obus[temp_w*0 +:temp_w];
assign v1068ibus[data_w*0 +:data_w] = c96obus[data_w*4 +:data_w];
assign c96ibus[temp_w*5 +:temp_w] = v1248obus[temp_w*1 +:temp_w];
assign v1248ibus[data_w*1 +:data_w] = c96obus[data_w*5 +:data_w];
assign c96ibus[temp_w*6 +:temp_w] = v1344obus[temp_w*0 +:temp_w];
assign v1344ibus[data_w*0 +:data_w] = c96obus[data_w*6 +:data_w];
assign c97ibus[temp_w*0 +:temp_w] = v124obus[temp_w*1 +:temp_w];
assign v124ibus[data_w*1 +:data_w] = c97obus[data_w*0 +:data_w];
assign c97ibus[temp_w*1 +:temp_w] = v503obus[temp_w*0 +:temp_w];
assign v503ibus[data_w*0 +:data_w] = c97obus[data_w*1 +:data_w];
assign c97ibus[temp_w*2 +:temp_w] = v656obus[temp_w*0 +:temp_w];
assign v656ibus[data_w*0 +:data_w] = c97obus[data_w*2 +:data_w];
assign c97ibus[temp_w*3 +:temp_w] = v682obus[temp_w*0 +:temp_w];
assign v682ibus[data_w*0 +:data_w] = c97obus[data_w*3 +:data_w];
assign c97ibus[temp_w*4 +:temp_w] = v1069obus[temp_w*0 +:temp_w];
assign v1069ibus[data_w*0 +:data_w] = c97obus[data_w*4 +:data_w];
assign c97ibus[temp_w*5 +:temp_w] = v1249obus[temp_w*1 +:temp_w];
assign v1249ibus[data_w*1 +:data_w] = c97obus[data_w*5 +:data_w];
assign c97ibus[temp_w*6 +:temp_w] = v1345obus[temp_w*0 +:temp_w];
assign v1345ibus[data_w*0 +:data_w] = c97obus[data_w*6 +:data_w];
assign c98ibus[temp_w*0 +:temp_w] = v125obus[temp_w*1 +:temp_w];
assign v125ibus[data_w*1 +:data_w] = c98obus[data_w*0 +:data_w];
assign c98ibus[temp_w*1 +:temp_w] = v504obus[temp_w*0 +:temp_w];
assign v504ibus[data_w*0 +:data_w] = c98obus[data_w*1 +:data_w];
assign c98ibus[temp_w*2 +:temp_w] = v657obus[temp_w*0 +:temp_w];
assign v657ibus[data_w*0 +:data_w] = c98obus[data_w*2 +:data_w];
assign c98ibus[temp_w*3 +:temp_w] = v683obus[temp_w*0 +:temp_w];
assign v683ibus[data_w*0 +:data_w] = c98obus[data_w*3 +:data_w];
assign c98ibus[temp_w*4 +:temp_w] = v1070obus[temp_w*0 +:temp_w];
assign v1070ibus[data_w*0 +:data_w] = c98obus[data_w*4 +:data_w];
assign c98ibus[temp_w*5 +:temp_w] = v1250obus[temp_w*1 +:temp_w];
assign v1250ibus[data_w*1 +:data_w] = c98obus[data_w*5 +:data_w];
assign c98ibus[temp_w*6 +:temp_w] = v1346obus[temp_w*0 +:temp_w];
assign v1346ibus[data_w*0 +:data_w] = c98obus[data_w*6 +:data_w];
assign c99ibus[temp_w*0 +:temp_w] = v126obus[temp_w*1 +:temp_w];
assign v126ibus[data_w*1 +:data_w] = c99obus[data_w*0 +:data_w];
assign c99ibus[temp_w*1 +:temp_w] = v505obus[temp_w*0 +:temp_w];
assign v505ibus[data_w*0 +:data_w] = c99obus[data_w*1 +:data_w];
assign c99ibus[temp_w*2 +:temp_w] = v658obus[temp_w*0 +:temp_w];
assign v658ibus[data_w*0 +:data_w] = c99obus[data_w*2 +:data_w];
assign c99ibus[temp_w*3 +:temp_w] = v684obus[temp_w*0 +:temp_w];
assign v684ibus[data_w*0 +:data_w] = c99obus[data_w*3 +:data_w];
assign c99ibus[temp_w*4 +:temp_w] = v1071obus[temp_w*0 +:temp_w];
assign v1071ibus[data_w*0 +:data_w] = c99obus[data_w*4 +:data_w];
assign c99ibus[temp_w*5 +:temp_w] = v1251obus[temp_w*1 +:temp_w];
assign v1251ibus[data_w*1 +:data_w] = c99obus[data_w*5 +:data_w];
assign c99ibus[temp_w*6 +:temp_w] = v1347obus[temp_w*0 +:temp_w];
assign v1347ibus[data_w*0 +:data_w] = c99obus[data_w*6 +:data_w];
assign c100ibus[temp_w*0 +:temp_w] = v127obus[temp_w*1 +:temp_w];
assign v127ibus[data_w*1 +:data_w] = c100obus[data_w*0 +:data_w];
assign c100ibus[temp_w*1 +:temp_w] = v506obus[temp_w*0 +:temp_w];
assign v506ibus[data_w*0 +:data_w] = c100obus[data_w*1 +:data_w];
assign c100ibus[temp_w*2 +:temp_w] = v659obus[temp_w*0 +:temp_w];
assign v659ibus[data_w*0 +:data_w] = c100obus[data_w*2 +:data_w];
assign c100ibus[temp_w*3 +:temp_w] = v685obus[temp_w*0 +:temp_w];
assign v685ibus[data_w*0 +:data_w] = c100obus[data_w*3 +:data_w];
assign c100ibus[temp_w*4 +:temp_w] = v1072obus[temp_w*0 +:temp_w];
assign v1072ibus[data_w*0 +:data_w] = c100obus[data_w*4 +:data_w];
assign c100ibus[temp_w*5 +:temp_w] = v1252obus[temp_w*1 +:temp_w];
assign v1252ibus[data_w*1 +:data_w] = c100obus[data_w*5 +:data_w];
assign c100ibus[temp_w*6 +:temp_w] = v1348obus[temp_w*0 +:temp_w];
assign v1348ibus[data_w*0 +:data_w] = c100obus[data_w*6 +:data_w];
assign c101ibus[temp_w*0 +:temp_w] = v128obus[temp_w*1 +:temp_w];
assign v128ibus[data_w*1 +:data_w] = c101obus[data_w*0 +:data_w];
assign c101ibus[temp_w*1 +:temp_w] = v507obus[temp_w*0 +:temp_w];
assign v507ibus[data_w*0 +:data_w] = c101obus[data_w*1 +:data_w];
assign c101ibus[temp_w*2 +:temp_w] = v660obus[temp_w*0 +:temp_w];
assign v660ibus[data_w*0 +:data_w] = c101obus[data_w*2 +:data_w];
assign c101ibus[temp_w*3 +:temp_w] = v686obus[temp_w*0 +:temp_w];
assign v686ibus[data_w*0 +:data_w] = c101obus[data_w*3 +:data_w];
assign c101ibus[temp_w*4 +:temp_w] = v1073obus[temp_w*0 +:temp_w];
assign v1073ibus[data_w*0 +:data_w] = c101obus[data_w*4 +:data_w];
assign c101ibus[temp_w*5 +:temp_w] = v1253obus[temp_w*1 +:temp_w];
assign v1253ibus[data_w*1 +:data_w] = c101obus[data_w*5 +:data_w];
assign c101ibus[temp_w*6 +:temp_w] = v1349obus[temp_w*0 +:temp_w];
assign v1349ibus[data_w*0 +:data_w] = c101obus[data_w*6 +:data_w];
assign c102ibus[temp_w*0 +:temp_w] = v129obus[temp_w*1 +:temp_w];
assign v129ibus[data_w*1 +:data_w] = c102obus[data_w*0 +:data_w];
assign c102ibus[temp_w*1 +:temp_w] = v508obus[temp_w*0 +:temp_w];
assign v508ibus[data_w*0 +:data_w] = c102obus[data_w*1 +:data_w];
assign c102ibus[temp_w*2 +:temp_w] = v661obus[temp_w*0 +:temp_w];
assign v661ibus[data_w*0 +:data_w] = c102obus[data_w*2 +:data_w];
assign c102ibus[temp_w*3 +:temp_w] = v687obus[temp_w*0 +:temp_w];
assign v687ibus[data_w*0 +:data_w] = c102obus[data_w*3 +:data_w];
assign c102ibus[temp_w*4 +:temp_w] = v1074obus[temp_w*0 +:temp_w];
assign v1074ibus[data_w*0 +:data_w] = c102obus[data_w*4 +:data_w];
assign c102ibus[temp_w*5 +:temp_w] = v1254obus[temp_w*1 +:temp_w];
assign v1254ibus[data_w*1 +:data_w] = c102obus[data_w*5 +:data_w];
assign c102ibus[temp_w*6 +:temp_w] = v1350obus[temp_w*0 +:temp_w];
assign v1350ibus[data_w*0 +:data_w] = c102obus[data_w*6 +:data_w];
assign c103ibus[temp_w*0 +:temp_w] = v130obus[temp_w*1 +:temp_w];
assign v130ibus[data_w*1 +:data_w] = c103obus[data_w*0 +:data_w];
assign c103ibus[temp_w*1 +:temp_w] = v509obus[temp_w*0 +:temp_w];
assign v509ibus[data_w*0 +:data_w] = c103obus[data_w*1 +:data_w];
assign c103ibus[temp_w*2 +:temp_w] = v662obus[temp_w*0 +:temp_w];
assign v662ibus[data_w*0 +:data_w] = c103obus[data_w*2 +:data_w];
assign c103ibus[temp_w*3 +:temp_w] = v688obus[temp_w*0 +:temp_w];
assign v688ibus[data_w*0 +:data_w] = c103obus[data_w*3 +:data_w];
assign c103ibus[temp_w*4 +:temp_w] = v1075obus[temp_w*0 +:temp_w];
assign v1075ibus[data_w*0 +:data_w] = c103obus[data_w*4 +:data_w];
assign c103ibus[temp_w*5 +:temp_w] = v1255obus[temp_w*1 +:temp_w];
assign v1255ibus[data_w*1 +:data_w] = c103obus[data_w*5 +:data_w];
assign c103ibus[temp_w*6 +:temp_w] = v1351obus[temp_w*0 +:temp_w];
assign v1351ibus[data_w*0 +:data_w] = c103obus[data_w*6 +:data_w];
assign c104ibus[temp_w*0 +:temp_w] = v131obus[temp_w*1 +:temp_w];
assign v131ibus[data_w*1 +:data_w] = c104obus[data_w*0 +:data_w];
assign c104ibus[temp_w*1 +:temp_w] = v510obus[temp_w*0 +:temp_w];
assign v510ibus[data_w*0 +:data_w] = c104obus[data_w*1 +:data_w];
assign c104ibus[temp_w*2 +:temp_w] = v663obus[temp_w*0 +:temp_w];
assign v663ibus[data_w*0 +:data_w] = c104obus[data_w*2 +:data_w];
assign c104ibus[temp_w*3 +:temp_w] = v689obus[temp_w*0 +:temp_w];
assign v689ibus[data_w*0 +:data_w] = c104obus[data_w*3 +:data_w];
assign c104ibus[temp_w*4 +:temp_w] = v1076obus[temp_w*0 +:temp_w];
assign v1076ibus[data_w*0 +:data_w] = c104obus[data_w*4 +:data_w];
assign c104ibus[temp_w*5 +:temp_w] = v1256obus[temp_w*1 +:temp_w];
assign v1256ibus[data_w*1 +:data_w] = c104obus[data_w*5 +:data_w];
assign c104ibus[temp_w*6 +:temp_w] = v1352obus[temp_w*0 +:temp_w];
assign v1352ibus[data_w*0 +:data_w] = c104obus[data_w*6 +:data_w];
assign c105ibus[temp_w*0 +:temp_w] = v132obus[temp_w*1 +:temp_w];
assign v132ibus[data_w*1 +:data_w] = c105obus[data_w*0 +:data_w];
assign c105ibus[temp_w*1 +:temp_w] = v511obus[temp_w*0 +:temp_w];
assign v511ibus[data_w*0 +:data_w] = c105obus[data_w*1 +:data_w];
assign c105ibus[temp_w*2 +:temp_w] = v664obus[temp_w*0 +:temp_w];
assign v664ibus[data_w*0 +:data_w] = c105obus[data_w*2 +:data_w];
assign c105ibus[temp_w*3 +:temp_w] = v690obus[temp_w*0 +:temp_w];
assign v690ibus[data_w*0 +:data_w] = c105obus[data_w*3 +:data_w];
assign c105ibus[temp_w*4 +:temp_w] = v1077obus[temp_w*0 +:temp_w];
assign v1077ibus[data_w*0 +:data_w] = c105obus[data_w*4 +:data_w];
assign c105ibus[temp_w*5 +:temp_w] = v1257obus[temp_w*1 +:temp_w];
assign v1257ibus[data_w*1 +:data_w] = c105obus[data_w*5 +:data_w];
assign c105ibus[temp_w*6 +:temp_w] = v1353obus[temp_w*0 +:temp_w];
assign v1353ibus[data_w*0 +:data_w] = c105obus[data_w*6 +:data_w];
assign c106ibus[temp_w*0 +:temp_w] = v133obus[temp_w*1 +:temp_w];
assign v133ibus[data_w*1 +:data_w] = c106obus[data_w*0 +:data_w];
assign c106ibus[temp_w*1 +:temp_w] = v512obus[temp_w*0 +:temp_w];
assign v512ibus[data_w*0 +:data_w] = c106obus[data_w*1 +:data_w];
assign c106ibus[temp_w*2 +:temp_w] = v665obus[temp_w*0 +:temp_w];
assign v665ibus[data_w*0 +:data_w] = c106obus[data_w*2 +:data_w];
assign c106ibus[temp_w*3 +:temp_w] = v691obus[temp_w*0 +:temp_w];
assign v691ibus[data_w*0 +:data_w] = c106obus[data_w*3 +:data_w];
assign c106ibus[temp_w*4 +:temp_w] = v1078obus[temp_w*0 +:temp_w];
assign v1078ibus[data_w*0 +:data_w] = c106obus[data_w*4 +:data_w];
assign c106ibus[temp_w*5 +:temp_w] = v1258obus[temp_w*1 +:temp_w];
assign v1258ibus[data_w*1 +:data_w] = c106obus[data_w*5 +:data_w];
assign c106ibus[temp_w*6 +:temp_w] = v1354obus[temp_w*0 +:temp_w];
assign v1354ibus[data_w*0 +:data_w] = c106obus[data_w*6 +:data_w];
assign c107ibus[temp_w*0 +:temp_w] = v134obus[temp_w*1 +:temp_w];
assign v134ibus[data_w*1 +:data_w] = c107obus[data_w*0 +:data_w];
assign c107ibus[temp_w*1 +:temp_w] = v513obus[temp_w*0 +:temp_w];
assign v513ibus[data_w*0 +:data_w] = c107obus[data_w*1 +:data_w];
assign c107ibus[temp_w*2 +:temp_w] = v666obus[temp_w*0 +:temp_w];
assign v666ibus[data_w*0 +:data_w] = c107obus[data_w*2 +:data_w];
assign c107ibus[temp_w*3 +:temp_w] = v692obus[temp_w*0 +:temp_w];
assign v692ibus[data_w*0 +:data_w] = c107obus[data_w*3 +:data_w];
assign c107ibus[temp_w*4 +:temp_w] = v1079obus[temp_w*0 +:temp_w];
assign v1079ibus[data_w*0 +:data_w] = c107obus[data_w*4 +:data_w];
assign c107ibus[temp_w*5 +:temp_w] = v1259obus[temp_w*1 +:temp_w];
assign v1259ibus[data_w*1 +:data_w] = c107obus[data_w*5 +:data_w];
assign c107ibus[temp_w*6 +:temp_w] = v1355obus[temp_w*0 +:temp_w];
assign v1355ibus[data_w*0 +:data_w] = c107obus[data_w*6 +:data_w];
assign c108ibus[temp_w*0 +:temp_w] = v135obus[temp_w*1 +:temp_w];
assign v135ibus[data_w*1 +:data_w] = c108obus[data_w*0 +:data_w];
assign c108ibus[temp_w*1 +:temp_w] = v514obus[temp_w*0 +:temp_w];
assign v514ibus[data_w*0 +:data_w] = c108obus[data_w*1 +:data_w];
assign c108ibus[temp_w*2 +:temp_w] = v667obus[temp_w*0 +:temp_w];
assign v667ibus[data_w*0 +:data_w] = c108obus[data_w*2 +:data_w];
assign c108ibus[temp_w*3 +:temp_w] = v693obus[temp_w*0 +:temp_w];
assign v693ibus[data_w*0 +:data_w] = c108obus[data_w*3 +:data_w];
assign c108ibus[temp_w*4 +:temp_w] = v1080obus[temp_w*0 +:temp_w];
assign v1080ibus[data_w*0 +:data_w] = c108obus[data_w*4 +:data_w];
assign c108ibus[temp_w*5 +:temp_w] = v1260obus[temp_w*1 +:temp_w];
assign v1260ibus[data_w*1 +:data_w] = c108obus[data_w*5 +:data_w];
assign c108ibus[temp_w*6 +:temp_w] = v1356obus[temp_w*0 +:temp_w];
assign v1356ibus[data_w*0 +:data_w] = c108obus[data_w*6 +:data_w];
assign c109ibus[temp_w*0 +:temp_w] = v136obus[temp_w*1 +:temp_w];
assign v136ibus[data_w*1 +:data_w] = c109obus[data_w*0 +:data_w];
assign c109ibus[temp_w*1 +:temp_w] = v515obus[temp_w*0 +:temp_w];
assign v515ibus[data_w*0 +:data_w] = c109obus[data_w*1 +:data_w];
assign c109ibus[temp_w*2 +:temp_w] = v668obus[temp_w*0 +:temp_w];
assign v668ibus[data_w*0 +:data_w] = c109obus[data_w*2 +:data_w];
assign c109ibus[temp_w*3 +:temp_w] = v694obus[temp_w*0 +:temp_w];
assign v694ibus[data_w*0 +:data_w] = c109obus[data_w*3 +:data_w];
assign c109ibus[temp_w*4 +:temp_w] = v1081obus[temp_w*0 +:temp_w];
assign v1081ibus[data_w*0 +:data_w] = c109obus[data_w*4 +:data_w];
assign c109ibus[temp_w*5 +:temp_w] = v1261obus[temp_w*1 +:temp_w];
assign v1261ibus[data_w*1 +:data_w] = c109obus[data_w*5 +:data_w];
assign c109ibus[temp_w*6 +:temp_w] = v1357obus[temp_w*0 +:temp_w];
assign v1357ibus[data_w*0 +:data_w] = c109obus[data_w*6 +:data_w];
assign c110ibus[temp_w*0 +:temp_w] = v137obus[temp_w*1 +:temp_w];
assign v137ibus[data_w*1 +:data_w] = c110obus[data_w*0 +:data_w];
assign c110ibus[temp_w*1 +:temp_w] = v516obus[temp_w*0 +:temp_w];
assign v516ibus[data_w*0 +:data_w] = c110obus[data_w*1 +:data_w];
assign c110ibus[temp_w*2 +:temp_w] = v669obus[temp_w*0 +:temp_w];
assign v669ibus[data_w*0 +:data_w] = c110obus[data_w*2 +:data_w];
assign c110ibus[temp_w*3 +:temp_w] = v695obus[temp_w*0 +:temp_w];
assign v695ibus[data_w*0 +:data_w] = c110obus[data_w*3 +:data_w];
assign c110ibus[temp_w*4 +:temp_w] = v1082obus[temp_w*0 +:temp_w];
assign v1082ibus[data_w*0 +:data_w] = c110obus[data_w*4 +:data_w];
assign c110ibus[temp_w*5 +:temp_w] = v1262obus[temp_w*1 +:temp_w];
assign v1262ibus[data_w*1 +:data_w] = c110obus[data_w*5 +:data_w];
assign c110ibus[temp_w*6 +:temp_w] = v1358obus[temp_w*0 +:temp_w];
assign v1358ibus[data_w*0 +:data_w] = c110obus[data_w*6 +:data_w];
assign c111ibus[temp_w*0 +:temp_w] = v138obus[temp_w*1 +:temp_w];
assign v138ibus[data_w*1 +:data_w] = c111obus[data_w*0 +:data_w];
assign c111ibus[temp_w*1 +:temp_w] = v517obus[temp_w*0 +:temp_w];
assign v517ibus[data_w*0 +:data_w] = c111obus[data_w*1 +:data_w];
assign c111ibus[temp_w*2 +:temp_w] = v670obus[temp_w*0 +:temp_w];
assign v670ibus[data_w*0 +:data_w] = c111obus[data_w*2 +:data_w];
assign c111ibus[temp_w*3 +:temp_w] = v696obus[temp_w*0 +:temp_w];
assign v696ibus[data_w*0 +:data_w] = c111obus[data_w*3 +:data_w];
assign c111ibus[temp_w*4 +:temp_w] = v1083obus[temp_w*0 +:temp_w];
assign v1083ibus[data_w*0 +:data_w] = c111obus[data_w*4 +:data_w];
assign c111ibus[temp_w*5 +:temp_w] = v1263obus[temp_w*1 +:temp_w];
assign v1263ibus[data_w*1 +:data_w] = c111obus[data_w*5 +:data_w];
assign c111ibus[temp_w*6 +:temp_w] = v1359obus[temp_w*0 +:temp_w];
assign v1359ibus[data_w*0 +:data_w] = c111obus[data_w*6 +:data_w];
assign c112ibus[temp_w*0 +:temp_w] = v139obus[temp_w*1 +:temp_w];
assign v139ibus[data_w*1 +:data_w] = c112obus[data_w*0 +:data_w];
assign c112ibus[temp_w*1 +:temp_w] = v518obus[temp_w*0 +:temp_w];
assign v518ibus[data_w*0 +:data_w] = c112obus[data_w*1 +:data_w];
assign c112ibus[temp_w*2 +:temp_w] = v671obus[temp_w*0 +:temp_w];
assign v671ibus[data_w*0 +:data_w] = c112obus[data_w*2 +:data_w];
assign c112ibus[temp_w*3 +:temp_w] = v697obus[temp_w*0 +:temp_w];
assign v697ibus[data_w*0 +:data_w] = c112obus[data_w*3 +:data_w];
assign c112ibus[temp_w*4 +:temp_w] = v1084obus[temp_w*0 +:temp_w];
assign v1084ibus[data_w*0 +:data_w] = c112obus[data_w*4 +:data_w];
assign c112ibus[temp_w*5 +:temp_w] = v1264obus[temp_w*1 +:temp_w];
assign v1264ibus[data_w*1 +:data_w] = c112obus[data_w*5 +:data_w];
assign c112ibus[temp_w*6 +:temp_w] = v1360obus[temp_w*0 +:temp_w];
assign v1360ibus[data_w*0 +:data_w] = c112obus[data_w*6 +:data_w];
assign c113ibus[temp_w*0 +:temp_w] = v140obus[temp_w*1 +:temp_w];
assign v140ibus[data_w*1 +:data_w] = c113obus[data_w*0 +:data_w];
assign c113ibus[temp_w*1 +:temp_w] = v519obus[temp_w*0 +:temp_w];
assign v519ibus[data_w*0 +:data_w] = c113obus[data_w*1 +:data_w];
assign c113ibus[temp_w*2 +:temp_w] = v576obus[temp_w*0 +:temp_w];
assign v576ibus[data_w*0 +:data_w] = c113obus[data_w*2 +:data_w];
assign c113ibus[temp_w*3 +:temp_w] = v698obus[temp_w*0 +:temp_w];
assign v698ibus[data_w*0 +:data_w] = c113obus[data_w*3 +:data_w];
assign c113ibus[temp_w*4 +:temp_w] = v1085obus[temp_w*0 +:temp_w];
assign v1085ibus[data_w*0 +:data_w] = c113obus[data_w*4 +:data_w];
assign c113ibus[temp_w*5 +:temp_w] = v1265obus[temp_w*1 +:temp_w];
assign v1265ibus[data_w*1 +:data_w] = c113obus[data_w*5 +:data_w];
assign c113ibus[temp_w*6 +:temp_w] = v1361obus[temp_w*0 +:temp_w];
assign v1361ibus[data_w*0 +:data_w] = c113obus[data_w*6 +:data_w];
assign c114ibus[temp_w*0 +:temp_w] = v141obus[temp_w*1 +:temp_w];
assign v141ibus[data_w*1 +:data_w] = c114obus[data_w*0 +:data_w];
assign c114ibus[temp_w*1 +:temp_w] = v520obus[temp_w*0 +:temp_w];
assign v520ibus[data_w*0 +:data_w] = c114obus[data_w*1 +:data_w];
assign c114ibus[temp_w*2 +:temp_w] = v577obus[temp_w*0 +:temp_w];
assign v577ibus[data_w*0 +:data_w] = c114obus[data_w*2 +:data_w];
assign c114ibus[temp_w*3 +:temp_w] = v699obus[temp_w*0 +:temp_w];
assign v699ibus[data_w*0 +:data_w] = c114obus[data_w*3 +:data_w];
assign c114ibus[temp_w*4 +:temp_w] = v1086obus[temp_w*0 +:temp_w];
assign v1086ibus[data_w*0 +:data_w] = c114obus[data_w*4 +:data_w];
assign c114ibus[temp_w*5 +:temp_w] = v1266obus[temp_w*1 +:temp_w];
assign v1266ibus[data_w*1 +:data_w] = c114obus[data_w*5 +:data_w];
assign c114ibus[temp_w*6 +:temp_w] = v1362obus[temp_w*0 +:temp_w];
assign v1362ibus[data_w*0 +:data_w] = c114obus[data_w*6 +:data_w];
assign c115ibus[temp_w*0 +:temp_w] = v142obus[temp_w*1 +:temp_w];
assign v142ibus[data_w*1 +:data_w] = c115obus[data_w*0 +:data_w];
assign c115ibus[temp_w*1 +:temp_w] = v521obus[temp_w*0 +:temp_w];
assign v521ibus[data_w*0 +:data_w] = c115obus[data_w*1 +:data_w];
assign c115ibus[temp_w*2 +:temp_w] = v578obus[temp_w*0 +:temp_w];
assign v578ibus[data_w*0 +:data_w] = c115obus[data_w*2 +:data_w];
assign c115ibus[temp_w*3 +:temp_w] = v700obus[temp_w*0 +:temp_w];
assign v700ibus[data_w*0 +:data_w] = c115obus[data_w*3 +:data_w];
assign c115ibus[temp_w*4 +:temp_w] = v1087obus[temp_w*0 +:temp_w];
assign v1087ibus[data_w*0 +:data_w] = c115obus[data_w*4 +:data_w];
assign c115ibus[temp_w*5 +:temp_w] = v1267obus[temp_w*1 +:temp_w];
assign v1267ibus[data_w*1 +:data_w] = c115obus[data_w*5 +:data_w];
assign c115ibus[temp_w*6 +:temp_w] = v1363obus[temp_w*0 +:temp_w];
assign v1363ibus[data_w*0 +:data_w] = c115obus[data_w*6 +:data_w];
assign c116ibus[temp_w*0 +:temp_w] = v143obus[temp_w*1 +:temp_w];
assign v143ibus[data_w*1 +:data_w] = c116obus[data_w*0 +:data_w];
assign c116ibus[temp_w*1 +:temp_w] = v522obus[temp_w*0 +:temp_w];
assign v522ibus[data_w*0 +:data_w] = c116obus[data_w*1 +:data_w];
assign c116ibus[temp_w*2 +:temp_w] = v579obus[temp_w*0 +:temp_w];
assign v579ibus[data_w*0 +:data_w] = c116obus[data_w*2 +:data_w];
assign c116ibus[temp_w*3 +:temp_w] = v701obus[temp_w*0 +:temp_w];
assign v701ibus[data_w*0 +:data_w] = c116obus[data_w*3 +:data_w];
assign c116ibus[temp_w*4 +:temp_w] = v1088obus[temp_w*0 +:temp_w];
assign v1088ibus[data_w*0 +:data_w] = c116obus[data_w*4 +:data_w];
assign c116ibus[temp_w*5 +:temp_w] = v1268obus[temp_w*1 +:temp_w];
assign v1268ibus[data_w*1 +:data_w] = c116obus[data_w*5 +:data_w];
assign c116ibus[temp_w*6 +:temp_w] = v1364obus[temp_w*0 +:temp_w];
assign v1364ibus[data_w*0 +:data_w] = c116obus[data_w*6 +:data_w];
assign c117ibus[temp_w*0 +:temp_w] = v144obus[temp_w*1 +:temp_w];
assign v144ibus[data_w*1 +:data_w] = c117obus[data_w*0 +:data_w];
assign c117ibus[temp_w*1 +:temp_w] = v523obus[temp_w*0 +:temp_w];
assign v523ibus[data_w*0 +:data_w] = c117obus[data_w*1 +:data_w];
assign c117ibus[temp_w*2 +:temp_w] = v580obus[temp_w*0 +:temp_w];
assign v580ibus[data_w*0 +:data_w] = c117obus[data_w*2 +:data_w];
assign c117ibus[temp_w*3 +:temp_w] = v702obus[temp_w*0 +:temp_w];
assign v702ibus[data_w*0 +:data_w] = c117obus[data_w*3 +:data_w];
assign c117ibus[temp_w*4 +:temp_w] = v1089obus[temp_w*0 +:temp_w];
assign v1089ibus[data_w*0 +:data_w] = c117obus[data_w*4 +:data_w];
assign c117ibus[temp_w*5 +:temp_w] = v1269obus[temp_w*1 +:temp_w];
assign v1269ibus[data_w*1 +:data_w] = c117obus[data_w*5 +:data_w];
assign c117ibus[temp_w*6 +:temp_w] = v1365obus[temp_w*0 +:temp_w];
assign v1365ibus[data_w*0 +:data_w] = c117obus[data_w*6 +:data_w];
assign c118ibus[temp_w*0 +:temp_w] = v145obus[temp_w*1 +:temp_w];
assign v145ibus[data_w*1 +:data_w] = c118obus[data_w*0 +:data_w];
assign c118ibus[temp_w*1 +:temp_w] = v524obus[temp_w*0 +:temp_w];
assign v524ibus[data_w*0 +:data_w] = c118obus[data_w*1 +:data_w];
assign c118ibus[temp_w*2 +:temp_w] = v581obus[temp_w*0 +:temp_w];
assign v581ibus[data_w*0 +:data_w] = c118obus[data_w*2 +:data_w];
assign c118ibus[temp_w*3 +:temp_w] = v703obus[temp_w*0 +:temp_w];
assign v703ibus[data_w*0 +:data_w] = c118obus[data_w*3 +:data_w];
assign c118ibus[temp_w*4 +:temp_w] = v1090obus[temp_w*0 +:temp_w];
assign v1090ibus[data_w*0 +:data_w] = c118obus[data_w*4 +:data_w];
assign c118ibus[temp_w*5 +:temp_w] = v1270obus[temp_w*1 +:temp_w];
assign v1270ibus[data_w*1 +:data_w] = c118obus[data_w*5 +:data_w];
assign c118ibus[temp_w*6 +:temp_w] = v1366obus[temp_w*0 +:temp_w];
assign v1366ibus[data_w*0 +:data_w] = c118obus[data_w*6 +:data_w];
assign c119ibus[temp_w*0 +:temp_w] = v146obus[temp_w*1 +:temp_w];
assign v146ibus[data_w*1 +:data_w] = c119obus[data_w*0 +:data_w];
assign c119ibus[temp_w*1 +:temp_w] = v525obus[temp_w*0 +:temp_w];
assign v525ibus[data_w*0 +:data_w] = c119obus[data_w*1 +:data_w];
assign c119ibus[temp_w*2 +:temp_w] = v582obus[temp_w*0 +:temp_w];
assign v582ibus[data_w*0 +:data_w] = c119obus[data_w*2 +:data_w];
assign c119ibus[temp_w*3 +:temp_w] = v704obus[temp_w*0 +:temp_w];
assign v704ibus[data_w*0 +:data_w] = c119obus[data_w*3 +:data_w];
assign c119ibus[temp_w*4 +:temp_w] = v1091obus[temp_w*0 +:temp_w];
assign v1091ibus[data_w*0 +:data_w] = c119obus[data_w*4 +:data_w];
assign c119ibus[temp_w*5 +:temp_w] = v1271obus[temp_w*1 +:temp_w];
assign v1271ibus[data_w*1 +:data_w] = c119obus[data_w*5 +:data_w];
assign c119ibus[temp_w*6 +:temp_w] = v1367obus[temp_w*0 +:temp_w];
assign v1367ibus[data_w*0 +:data_w] = c119obus[data_w*6 +:data_w];
assign c120ibus[temp_w*0 +:temp_w] = v147obus[temp_w*1 +:temp_w];
assign v147ibus[data_w*1 +:data_w] = c120obus[data_w*0 +:data_w];
assign c120ibus[temp_w*1 +:temp_w] = v526obus[temp_w*0 +:temp_w];
assign v526ibus[data_w*0 +:data_w] = c120obus[data_w*1 +:data_w];
assign c120ibus[temp_w*2 +:temp_w] = v583obus[temp_w*0 +:temp_w];
assign v583ibus[data_w*0 +:data_w] = c120obus[data_w*2 +:data_w];
assign c120ibus[temp_w*3 +:temp_w] = v705obus[temp_w*0 +:temp_w];
assign v705ibus[data_w*0 +:data_w] = c120obus[data_w*3 +:data_w];
assign c120ibus[temp_w*4 +:temp_w] = v1092obus[temp_w*0 +:temp_w];
assign v1092ibus[data_w*0 +:data_w] = c120obus[data_w*4 +:data_w];
assign c120ibus[temp_w*5 +:temp_w] = v1272obus[temp_w*1 +:temp_w];
assign v1272ibus[data_w*1 +:data_w] = c120obus[data_w*5 +:data_w];
assign c120ibus[temp_w*6 +:temp_w] = v1368obus[temp_w*0 +:temp_w];
assign v1368ibus[data_w*0 +:data_w] = c120obus[data_w*6 +:data_w];
assign c121ibus[temp_w*0 +:temp_w] = v148obus[temp_w*1 +:temp_w];
assign v148ibus[data_w*1 +:data_w] = c121obus[data_w*0 +:data_w];
assign c121ibus[temp_w*1 +:temp_w] = v527obus[temp_w*0 +:temp_w];
assign v527ibus[data_w*0 +:data_w] = c121obus[data_w*1 +:data_w];
assign c121ibus[temp_w*2 +:temp_w] = v584obus[temp_w*0 +:temp_w];
assign v584ibus[data_w*0 +:data_w] = c121obus[data_w*2 +:data_w];
assign c121ibus[temp_w*3 +:temp_w] = v706obus[temp_w*0 +:temp_w];
assign v706ibus[data_w*0 +:data_w] = c121obus[data_w*3 +:data_w];
assign c121ibus[temp_w*4 +:temp_w] = v1093obus[temp_w*0 +:temp_w];
assign v1093ibus[data_w*0 +:data_w] = c121obus[data_w*4 +:data_w];
assign c121ibus[temp_w*5 +:temp_w] = v1273obus[temp_w*1 +:temp_w];
assign v1273ibus[data_w*1 +:data_w] = c121obus[data_w*5 +:data_w];
assign c121ibus[temp_w*6 +:temp_w] = v1369obus[temp_w*0 +:temp_w];
assign v1369ibus[data_w*0 +:data_w] = c121obus[data_w*6 +:data_w];
assign c122ibus[temp_w*0 +:temp_w] = v149obus[temp_w*1 +:temp_w];
assign v149ibus[data_w*1 +:data_w] = c122obus[data_w*0 +:data_w];
assign c122ibus[temp_w*1 +:temp_w] = v528obus[temp_w*0 +:temp_w];
assign v528ibus[data_w*0 +:data_w] = c122obus[data_w*1 +:data_w];
assign c122ibus[temp_w*2 +:temp_w] = v585obus[temp_w*0 +:temp_w];
assign v585ibus[data_w*0 +:data_w] = c122obus[data_w*2 +:data_w];
assign c122ibus[temp_w*3 +:temp_w] = v707obus[temp_w*0 +:temp_w];
assign v707ibus[data_w*0 +:data_w] = c122obus[data_w*3 +:data_w];
assign c122ibus[temp_w*4 +:temp_w] = v1094obus[temp_w*0 +:temp_w];
assign v1094ibus[data_w*0 +:data_w] = c122obus[data_w*4 +:data_w];
assign c122ibus[temp_w*5 +:temp_w] = v1274obus[temp_w*1 +:temp_w];
assign v1274ibus[data_w*1 +:data_w] = c122obus[data_w*5 +:data_w];
assign c122ibus[temp_w*6 +:temp_w] = v1370obus[temp_w*0 +:temp_w];
assign v1370ibus[data_w*0 +:data_w] = c122obus[data_w*6 +:data_w];
assign c123ibus[temp_w*0 +:temp_w] = v150obus[temp_w*1 +:temp_w];
assign v150ibus[data_w*1 +:data_w] = c123obus[data_w*0 +:data_w];
assign c123ibus[temp_w*1 +:temp_w] = v529obus[temp_w*0 +:temp_w];
assign v529ibus[data_w*0 +:data_w] = c123obus[data_w*1 +:data_w];
assign c123ibus[temp_w*2 +:temp_w] = v586obus[temp_w*0 +:temp_w];
assign v586ibus[data_w*0 +:data_w] = c123obus[data_w*2 +:data_w];
assign c123ibus[temp_w*3 +:temp_w] = v708obus[temp_w*0 +:temp_w];
assign v708ibus[data_w*0 +:data_w] = c123obus[data_w*3 +:data_w];
assign c123ibus[temp_w*4 +:temp_w] = v1095obus[temp_w*0 +:temp_w];
assign v1095ibus[data_w*0 +:data_w] = c123obus[data_w*4 +:data_w];
assign c123ibus[temp_w*5 +:temp_w] = v1275obus[temp_w*1 +:temp_w];
assign v1275ibus[data_w*1 +:data_w] = c123obus[data_w*5 +:data_w];
assign c123ibus[temp_w*6 +:temp_w] = v1371obus[temp_w*0 +:temp_w];
assign v1371ibus[data_w*0 +:data_w] = c123obus[data_w*6 +:data_w];
assign c124ibus[temp_w*0 +:temp_w] = v151obus[temp_w*1 +:temp_w];
assign v151ibus[data_w*1 +:data_w] = c124obus[data_w*0 +:data_w];
assign c124ibus[temp_w*1 +:temp_w] = v530obus[temp_w*0 +:temp_w];
assign v530ibus[data_w*0 +:data_w] = c124obus[data_w*1 +:data_w];
assign c124ibus[temp_w*2 +:temp_w] = v587obus[temp_w*0 +:temp_w];
assign v587ibus[data_w*0 +:data_w] = c124obus[data_w*2 +:data_w];
assign c124ibus[temp_w*3 +:temp_w] = v709obus[temp_w*0 +:temp_w];
assign v709ibus[data_w*0 +:data_w] = c124obus[data_w*3 +:data_w];
assign c124ibus[temp_w*4 +:temp_w] = v1096obus[temp_w*0 +:temp_w];
assign v1096ibus[data_w*0 +:data_w] = c124obus[data_w*4 +:data_w];
assign c124ibus[temp_w*5 +:temp_w] = v1276obus[temp_w*1 +:temp_w];
assign v1276ibus[data_w*1 +:data_w] = c124obus[data_w*5 +:data_w];
assign c124ibus[temp_w*6 +:temp_w] = v1372obus[temp_w*0 +:temp_w];
assign v1372ibus[data_w*0 +:data_w] = c124obus[data_w*6 +:data_w];
assign c125ibus[temp_w*0 +:temp_w] = v152obus[temp_w*1 +:temp_w];
assign v152ibus[data_w*1 +:data_w] = c125obus[data_w*0 +:data_w];
assign c125ibus[temp_w*1 +:temp_w] = v531obus[temp_w*0 +:temp_w];
assign v531ibus[data_w*0 +:data_w] = c125obus[data_w*1 +:data_w];
assign c125ibus[temp_w*2 +:temp_w] = v588obus[temp_w*0 +:temp_w];
assign v588ibus[data_w*0 +:data_w] = c125obus[data_w*2 +:data_w];
assign c125ibus[temp_w*3 +:temp_w] = v710obus[temp_w*0 +:temp_w];
assign v710ibus[data_w*0 +:data_w] = c125obus[data_w*3 +:data_w];
assign c125ibus[temp_w*4 +:temp_w] = v1097obus[temp_w*0 +:temp_w];
assign v1097ibus[data_w*0 +:data_w] = c125obus[data_w*4 +:data_w];
assign c125ibus[temp_w*5 +:temp_w] = v1277obus[temp_w*1 +:temp_w];
assign v1277ibus[data_w*1 +:data_w] = c125obus[data_w*5 +:data_w];
assign c125ibus[temp_w*6 +:temp_w] = v1373obus[temp_w*0 +:temp_w];
assign v1373ibus[data_w*0 +:data_w] = c125obus[data_w*6 +:data_w];
assign c126ibus[temp_w*0 +:temp_w] = v153obus[temp_w*1 +:temp_w];
assign v153ibus[data_w*1 +:data_w] = c126obus[data_w*0 +:data_w];
assign c126ibus[temp_w*1 +:temp_w] = v532obus[temp_w*0 +:temp_w];
assign v532ibus[data_w*0 +:data_w] = c126obus[data_w*1 +:data_w];
assign c126ibus[temp_w*2 +:temp_w] = v589obus[temp_w*0 +:temp_w];
assign v589ibus[data_w*0 +:data_w] = c126obus[data_w*2 +:data_w];
assign c126ibus[temp_w*3 +:temp_w] = v711obus[temp_w*0 +:temp_w];
assign v711ibus[data_w*0 +:data_w] = c126obus[data_w*3 +:data_w];
assign c126ibus[temp_w*4 +:temp_w] = v1098obus[temp_w*0 +:temp_w];
assign v1098ibus[data_w*0 +:data_w] = c126obus[data_w*4 +:data_w];
assign c126ibus[temp_w*5 +:temp_w] = v1278obus[temp_w*1 +:temp_w];
assign v1278ibus[data_w*1 +:data_w] = c126obus[data_w*5 +:data_w];
assign c126ibus[temp_w*6 +:temp_w] = v1374obus[temp_w*0 +:temp_w];
assign v1374ibus[data_w*0 +:data_w] = c126obus[data_w*6 +:data_w];
assign c127ibus[temp_w*0 +:temp_w] = v154obus[temp_w*1 +:temp_w];
assign v154ibus[data_w*1 +:data_w] = c127obus[data_w*0 +:data_w];
assign c127ibus[temp_w*1 +:temp_w] = v533obus[temp_w*0 +:temp_w];
assign v533ibus[data_w*0 +:data_w] = c127obus[data_w*1 +:data_w];
assign c127ibus[temp_w*2 +:temp_w] = v590obus[temp_w*0 +:temp_w];
assign v590ibus[data_w*0 +:data_w] = c127obus[data_w*2 +:data_w];
assign c127ibus[temp_w*3 +:temp_w] = v712obus[temp_w*0 +:temp_w];
assign v712ibus[data_w*0 +:data_w] = c127obus[data_w*3 +:data_w];
assign c127ibus[temp_w*4 +:temp_w] = v1099obus[temp_w*0 +:temp_w];
assign v1099ibus[data_w*0 +:data_w] = c127obus[data_w*4 +:data_w];
assign c127ibus[temp_w*5 +:temp_w] = v1279obus[temp_w*1 +:temp_w];
assign v1279ibus[data_w*1 +:data_w] = c127obus[data_w*5 +:data_w];
assign c127ibus[temp_w*6 +:temp_w] = v1375obus[temp_w*0 +:temp_w];
assign v1375ibus[data_w*0 +:data_w] = c127obus[data_w*6 +:data_w];
assign c128ibus[temp_w*0 +:temp_w] = v155obus[temp_w*1 +:temp_w];
assign v155ibus[data_w*1 +:data_w] = c128obus[data_w*0 +:data_w];
assign c128ibus[temp_w*1 +:temp_w] = v534obus[temp_w*0 +:temp_w];
assign v534ibus[data_w*0 +:data_w] = c128obus[data_w*1 +:data_w];
assign c128ibus[temp_w*2 +:temp_w] = v591obus[temp_w*0 +:temp_w];
assign v591ibus[data_w*0 +:data_w] = c128obus[data_w*2 +:data_w];
assign c128ibus[temp_w*3 +:temp_w] = v713obus[temp_w*0 +:temp_w];
assign v713ibus[data_w*0 +:data_w] = c128obus[data_w*3 +:data_w];
assign c128ibus[temp_w*4 +:temp_w] = v1100obus[temp_w*0 +:temp_w];
assign v1100ibus[data_w*0 +:data_w] = c128obus[data_w*4 +:data_w];
assign c128ibus[temp_w*5 +:temp_w] = v1280obus[temp_w*1 +:temp_w];
assign v1280ibus[data_w*1 +:data_w] = c128obus[data_w*5 +:data_w];
assign c128ibus[temp_w*6 +:temp_w] = v1376obus[temp_w*0 +:temp_w];
assign v1376ibus[data_w*0 +:data_w] = c128obus[data_w*6 +:data_w];
assign c129ibus[temp_w*0 +:temp_w] = v156obus[temp_w*1 +:temp_w];
assign v156ibus[data_w*1 +:data_w] = c129obus[data_w*0 +:data_w];
assign c129ibus[temp_w*1 +:temp_w] = v535obus[temp_w*0 +:temp_w];
assign v535ibus[data_w*0 +:data_w] = c129obus[data_w*1 +:data_w];
assign c129ibus[temp_w*2 +:temp_w] = v592obus[temp_w*0 +:temp_w];
assign v592ibus[data_w*0 +:data_w] = c129obus[data_w*2 +:data_w];
assign c129ibus[temp_w*3 +:temp_w] = v714obus[temp_w*0 +:temp_w];
assign v714ibus[data_w*0 +:data_w] = c129obus[data_w*3 +:data_w];
assign c129ibus[temp_w*4 +:temp_w] = v1101obus[temp_w*0 +:temp_w];
assign v1101ibus[data_w*0 +:data_w] = c129obus[data_w*4 +:data_w];
assign c129ibus[temp_w*5 +:temp_w] = v1281obus[temp_w*1 +:temp_w];
assign v1281ibus[data_w*1 +:data_w] = c129obus[data_w*5 +:data_w];
assign c129ibus[temp_w*6 +:temp_w] = v1377obus[temp_w*0 +:temp_w];
assign v1377ibus[data_w*0 +:data_w] = c129obus[data_w*6 +:data_w];
assign c130ibus[temp_w*0 +:temp_w] = v157obus[temp_w*1 +:temp_w];
assign v157ibus[data_w*1 +:data_w] = c130obus[data_w*0 +:data_w];
assign c130ibus[temp_w*1 +:temp_w] = v536obus[temp_w*0 +:temp_w];
assign v536ibus[data_w*0 +:data_w] = c130obus[data_w*1 +:data_w];
assign c130ibus[temp_w*2 +:temp_w] = v593obus[temp_w*0 +:temp_w];
assign v593ibus[data_w*0 +:data_w] = c130obus[data_w*2 +:data_w];
assign c130ibus[temp_w*3 +:temp_w] = v715obus[temp_w*0 +:temp_w];
assign v715ibus[data_w*0 +:data_w] = c130obus[data_w*3 +:data_w];
assign c130ibus[temp_w*4 +:temp_w] = v1102obus[temp_w*0 +:temp_w];
assign v1102ibus[data_w*0 +:data_w] = c130obus[data_w*4 +:data_w];
assign c130ibus[temp_w*5 +:temp_w] = v1282obus[temp_w*1 +:temp_w];
assign v1282ibus[data_w*1 +:data_w] = c130obus[data_w*5 +:data_w];
assign c130ibus[temp_w*6 +:temp_w] = v1378obus[temp_w*0 +:temp_w];
assign v1378ibus[data_w*0 +:data_w] = c130obus[data_w*6 +:data_w];
assign c131ibus[temp_w*0 +:temp_w] = v158obus[temp_w*1 +:temp_w];
assign v158ibus[data_w*1 +:data_w] = c131obus[data_w*0 +:data_w];
assign c131ibus[temp_w*1 +:temp_w] = v537obus[temp_w*0 +:temp_w];
assign v537ibus[data_w*0 +:data_w] = c131obus[data_w*1 +:data_w];
assign c131ibus[temp_w*2 +:temp_w] = v594obus[temp_w*0 +:temp_w];
assign v594ibus[data_w*0 +:data_w] = c131obus[data_w*2 +:data_w];
assign c131ibus[temp_w*3 +:temp_w] = v716obus[temp_w*0 +:temp_w];
assign v716ibus[data_w*0 +:data_w] = c131obus[data_w*3 +:data_w];
assign c131ibus[temp_w*4 +:temp_w] = v1103obus[temp_w*0 +:temp_w];
assign v1103ibus[data_w*0 +:data_w] = c131obus[data_w*4 +:data_w];
assign c131ibus[temp_w*5 +:temp_w] = v1283obus[temp_w*1 +:temp_w];
assign v1283ibus[data_w*1 +:data_w] = c131obus[data_w*5 +:data_w];
assign c131ibus[temp_w*6 +:temp_w] = v1379obus[temp_w*0 +:temp_w];
assign v1379ibus[data_w*0 +:data_w] = c131obus[data_w*6 +:data_w];
assign c132ibus[temp_w*0 +:temp_w] = v159obus[temp_w*1 +:temp_w];
assign v159ibus[data_w*1 +:data_w] = c132obus[data_w*0 +:data_w];
assign c132ibus[temp_w*1 +:temp_w] = v538obus[temp_w*0 +:temp_w];
assign v538ibus[data_w*0 +:data_w] = c132obus[data_w*1 +:data_w];
assign c132ibus[temp_w*2 +:temp_w] = v595obus[temp_w*0 +:temp_w];
assign v595ibus[data_w*0 +:data_w] = c132obus[data_w*2 +:data_w];
assign c132ibus[temp_w*3 +:temp_w] = v717obus[temp_w*0 +:temp_w];
assign v717ibus[data_w*0 +:data_w] = c132obus[data_w*3 +:data_w];
assign c132ibus[temp_w*4 +:temp_w] = v1104obus[temp_w*0 +:temp_w];
assign v1104ibus[data_w*0 +:data_w] = c132obus[data_w*4 +:data_w];
assign c132ibus[temp_w*5 +:temp_w] = v1284obus[temp_w*1 +:temp_w];
assign v1284ibus[data_w*1 +:data_w] = c132obus[data_w*5 +:data_w];
assign c132ibus[temp_w*6 +:temp_w] = v1380obus[temp_w*0 +:temp_w];
assign v1380ibus[data_w*0 +:data_w] = c132obus[data_w*6 +:data_w];
assign c133ibus[temp_w*0 +:temp_w] = v160obus[temp_w*1 +:temp_w];
assign v160ibus[data_w*1 +:data_w] = c133obus[data_w*0 +:data_w];
assign c133ibus[temp_w*1 +:temp_w] = v539obus[temp_w*0 +:temp_w];
assign v539ibus[data_w*0 +:data_w] = c133obus[data_w*1 +:data_w];
assign c133ibus[temp_w*2 +:temp_w] = v596obus[temp_w*0 +:temp_w];
assign v596ibus[data_w*0 +:data_w] = c133obus[data_w*2 +:data_w];
assign c133ibus[temp_w*3 +:temp_w] = v718obus[temp_w*0 +:temp_w];
assign v718ibus[data_w*0 +:data_w] = c133obus[data_w*3 +:data_w];
assign c133ibus[temp_w*4 +:temp_w] = v1105obus[temp_w*0 +:temp_w];
assign v1105ibus[data_w*0 +:data_w] = c133obus[data_w*4 +:data_w];
assign c133ibus[temp_w*5 +:temp_w] = v1285obus[temp_w*1 +:temp_w];
assign v1285ibus[data_w*1 +:data_w] = c133obus[data_w*5 +:data_w];
assign c133ibus[temp_w*6 +:temp_w] = v1381obus[temp_w*0 +:temp_w];
assign v1381ibus[data_w*0 +:data_w] = c133obus[data_w*6 +:data_w];
assign c134ibus[temp_w*0 +:temp_w] = v161obus[temp_w*1 +:temp_w];
assign v161ibus[data_w*1 +:data_w] = c134obus[data_w*0 +:data_w];
assign c134ibus[temp_w*1 +:temp_w] = v540obus[temp_w*0 +:temp_w];
assign v540ibus[data_w*0 +:data_w] = c134obus[data_w*1 +:data_w];
assign c134ibus[temp_w*2 +:temp_w] = v597obus[temp_w*0 +:temp_w];
assign v597ibus[data_w*0 +:data_w] = c134obus[data_w*2 +:data_w];
assign c134ibus[temp_w*3 +:temp_w] = v719obus[temp_w*0 +:temp_w];
assign v719ibus[data_w*0 +:data_w] = c134obus[data_w*3 +:data_w];
assign c134ibus[temp_w*4 +:temp_w] = v1106obus[temp_w*0 +:temp_w];
assign v1106ibus[data_w*0 +:data_w] = c134obus[data_w*4 +:data_w];
assign c134ibus[temp_w*5 +:temp_w] = v1286obus[temp_w*1 +:temp_w];
assign v1286ibus[data_w*1 +:data_w] = c134obus[data_w*5 +:data_w];
assign c134ibus[temp_w*6 +:temp_w] = v1382obus[temp_w*0 +:temp_w];
assign v1382ibus[data_w*0 +:data_w] = c134obus[data_w*6 +:data_w];
assign c135ibus[temp_w*0 +:temp_w] = v162obus[temp_w*1 +:temp_w];
assign v162ibus[data_w*1 +:data_w] = c135obus[data_w*0 +:data_w];
assign c135ibus[temp_w*1 +:temp_w] = v541obus[temp_w*0 +:temp_w];
assign v541ibus[data_w*0 +:data_w] = c135obus[data_w*1 +:data_w];
assign c135ibus[temp_w*2 +:temp_w] = v598obus[temp_w*0 +:temp_w];
assign v598ibus[data_w*0 +:data_w] = c135obus[data_w*2 +:data_w];
assign c135ibus[temp_w*3 +:temp_w] = v720obus[temp_w*0 +:temp_w];
assign v720ibus[data_w*0 +:data_w] = c135obus[data_w*3 +:data_w];
assign c135ibus[temp_w*4 +:temp_w] = v1107obus[temp_w*0 +:temp_w];
assign v1107ibus[data_w*0 +:data_w] = c135obus[data_w*4 +:data_w];
assign c135ibus[temp_w*5 +:temp_w] = v1287obus[temp_w*1 +:temp_w];
assign v1287ibus[data_w*1 +:data_w] = c135obus[data_w*5 +:data_w];
assign c135ibus[temp_w*6 +:temp_w] = v1383obus[temp_w*0 +:temp_w];
assign v1383ibus[data_w*0 +:data_w] = c135obus[data_w*6 +:data_w];
assign c136ibus[temp_w*0 +:temp_w] = v163obus[temp_w*1 +:temp_w];
assign v163ibus[data_w*1 +:data_w] = c136obus[data_w*0 +:data_w];
assign c136ibus[temp_w*1 +:temp_w] = v542obus[temp_w*0 +:temp_w];
assign v542ibus[data_w*0 +:data_w] = c136obus[data_w*1 +:data_w];
assign c136ibus[temp_w*2 +:temp_w] = v599obus[temp_w*0 +:temp_w];
assign v599ibus[data_w*0 +:data_w] = c136obus[data_w*2 +:data_w];
assign c136ibus[temp_w*3 +:temp_w] = v721obus[temp_w*0 +:temp_w];
assign v721ibus[data_w*0 +:data_w] = c136obus[data_w*3 +:data_w];
assign c136ibus[temp_w*4 +:temp_w] = v1108obus[temp_w*0 +:temp_w];
assign v1108ibus[data_w*0 +:data_w] = c136obus[data_w*4 +:data_w];
assign c136ibus[temp_w*5 +:temp_w] = v1288obus[temp_w*1 +:temp_w];
assign v1288ibus[data_w*1 +:data_w] = c136obus[data_w*5 +:data_w];
assign c136ibus[temp_w*6 +:temp_w] = v1384obus[temp_w*0 +:temp_w];
assign v1384ibus[data_w*0 +:data_w] = c136obus[data_w*6 +:data_w];
assign c137ibus[temp_w*0 +:temp_w] = v164obus[temp_w*1 +:temp_w];
assign v164ibus[data_w*1 +:data_w] = c137obus[data_w*0 +:data_w];
assign c137ibus[temp_w*1 +:temp_w] = v543obus[temp_w*0 +:temp_w];
assign v543ibus[data_w*0 +:data_w] = c137obus[data_w*1 +:data_w];
assign c137ibus[temp_w*2 +:temp_w] = v600obus[temp_w*0 +:temp_w];
assign v600ibus[data_w*0 +:data_w] = c137obus[data_w*2 +:data_w];
assign c137ibus[temp_w*3 +:temp_w] = v722obus[temp_w*0 +:temp_w];
assign v722ibus[data_w*0 +:data_w] = c137obus[data_w*3 +:data_w];
assign c137ibus[temp_w*4 +:temp_w] = v1109obus[temp_w*0 +:temp_w];
assign v1109ibus[data_w*0 +:data_w] = c137obus[data_w*4 +:data_w];
assign c137ibus[temp_w*5 +:temp_w] = v1289obus[temp_w*1 +:temp_w];
assign v1289ibus[data_w*1 +:data_w] = c137obus[data_w*5 +:data_w];
assign c137ibus[temp_w*6 +:temp_w] = v1385obus[temp_w*0 +:temp_w];
assign v1385ibus[data_w*0 +:data_w] = c137obus[data_w*6 +:data_w];
assign c138ibus[temp_w*0 +:temp_w] = v165obus[temp_w*1 +:temp_w];
assign v165ibus[data_w*1 +:data_w] = c138obus[data_w*0 +:data_w];
assign c138ibus[temp_w*1 +:temp_w] = v544obus[temp_w*0 +:temp_w];
assign v544ibus[data_w*0 +:data_w] = c138obus[data_w*1 +:data_w];
assign c138ibus[temp_w*2 +:temp_w] = v601obus[temp_w*0 +:temp_w];
assign v601ibus[data_w*0 +:data_w] = c138obus[data_w*2 +:data_w];
assign c138ibus[temp_w*3 +:temp_w] = v723obus[temp_w*0 +:temp_w];
assign v723ibus[data_w*0 +:data_w] = c138obus[data_w*3 +:data_w];
assign c138ibus[temp_w*4 +:temp_w] = v1110obus[temp_w*0 +:temp_w];
assign v1110ibus[data_w*0 +:data_w] = c138obus[data_w*4 +:data_w];
assign c138ibus[temp_w*5 +:temp_w] = v1290obus[temp_w*1 +:temp_w];
assign v1290ibus[data_w*1 +:data_w] = c138obus[data_w*5 +:data_w];
assign c138ibus[temp_w*6 +:temp_w] = v1386obus[temp_w*0 +:temp_w];
assign v1386ibus[data_w*0 +:data_w] = c138obus[data_w*6 +:data_w];
assign c139ibus[temp_w*0 +:temp_w] = v166obus[temp_w*1 +:temp_w];
assign v166ibus[data_w*1 +:data_w] = c139obus[data_w*0 +:data_w];
assign c139ibus[temp_w*1 +:temp_w] = v545obus[temp_w*0 +:temp_w];
assign v545ibus[data_w*0 +:data_w] = c139obus[data_w*1 +:data_w];
assign c139ibus[temp_w*2 +:temp_w] = v602obus[temp_w*0 +:temp_w];
assign v602ibus[data_w*0 +:data_w] = c139obus[data_w*2 +:data_w];
assign c139ibus[temp_w*3 +:temp_w] = v724obus[temp_w*0 +:temp_w];
assign v724ibus[data_w*0 +:data_w] = c139obus[data_w*3 +:data_w];
assign c139ibus[temp_w*4 +:temp_w] = v1111obus[temp_w*0 +:temp_w];
assign v1111ibus[data_w*0 +:data_w] = c139obus[data_w*4 +:data_w];
assign c139ibus[temp_w*5 +:temp_w] = v1291obus[temp_w*1 +:temp_w];
assign v1291ibus[data_w*1 +:data_w] = c139obus[data_w*5 +:data_w];
assign c139ibus[temp_w*6 +:temp_w] = v1387obus[temp_w*0 +:temp_w];
assign v1387ibus[data_w*0 +:data_w] = c139obus[data_w*6 +:data_w];
assign c140ibus[temp_w*0 +:temp_w] = v167obus[temp_w*1 +:temp_w];
assign v167ibus[data_w*1 +:data_w] = c140obus[data_w*0 +:data_w];
assign c140ibus[temp_w*1 +:temp_w] = v546obus[temp_w*0 +:temp_w];
assign v546ibus[data_w*0 +:data_w] = c140obus[data_w*1 +:data_w];
assign c140ibus[temp_w*2 +:temp_w] = v603obus[temp_w*0 +:temp_w];
assign v603ibus[data_w*0 +:data_w] = c140obus[data_w*2 +:data_w];
assign c140ibus[temp_w*3 +:temp_w] = v725obus[temp_w*0 +:temp_w];
assign v725ibus[data_w*0 +:data_w] = c140obus[data_w*3 +:data_w];
assign c140ibus[temp_w*4 +:temp_w] = v1112obus[temp_w*0 +:temp_w];
assign v1112ibus[data_w*0 +:data_w] = c140obus[data_w*4 +:data_w];
assign c140ibus[temp_w*5 +:temp_w] = v1292obus[temp_w*1 +:temp_w];
assign v1292ibus[data_w*1 +:data_w] = c140obus[data_w*5 +:data_w];
assign c140ibus[temp_w*6 +:temp_w] = v1388obus[temp_w*0 +:temp_w];
assign v1388ibus[data_w*0 +:data_w] = c140obus[data_w*6 +:data_w];
assign c141ibus[temp_w*0 +:temp_w] = v168obus[temp_w*1 +:temp_w];
assign v168ibus[data_w*1 +:data_w] = c141obus[data_w*0 +:data_w];
assign c141ibus[temp_w*1 +:temp_w] = v547obus[temp_w*0 +:temp_w];
assign v547ibus[data_w*0 +:data_w] = c141obus[data_w*1 +:data_w];
assign c141ibus[temp_w*2 +:temp_w] = v604obus[temp_w*0 +:temp_w];
assign v604ibus[data_w*0 +:data_w] = c141obus[data_w*2 +:data_w];
assign c141ibus[temp_w*3 +:temp_w] = v726obus[temp_w*0 +:temp_w];
assign v726ibus[data_w*0 +:data_w] = c141obus[data_w*3 +:data_w];
assign c141ibus[temp_w*4 +:temp_w] = v1113obus[temp_w*0 +:temp_w];
assign v1113ibus[data_w*0 +:data_w] = c141obus[data_w*4 +:data_w];
assign c141ibus[temp_w*5 +:temp_w] = v1293obus[temp_w*1 +:temp_w];
assign v1293ibus[data_w*1 +:data_w] = c141obus[data_w*5 +:data_w];
assign c141ibus[temp_w*6 +:temp_w] = v1389obus[temp_w*0 +:temp_w];
assign v1389ibus[data_w*0 +:data_w] = c141obus[data_w*6 +:data_w];
assign c142ibus[temp_w*0 +:temp_w] = v169obus[temp_w*1 +:temp_w];
assign v169ibus[data_w*1 +:data_w] = c142obus[data_w*0 +:data_w];
assign c142ibus[temp_w*1 +:temp_w] = v548obus[temp_w*0 +:temp_w];
assign v548ibus[data_w*0 +:data_w] = c142obus[data_w*1 +:data_w];
assign c142ibus[temp_w*2 +:temp_w] = v605obus[temp_w*0 +:temp_w];
assign v605ibus[data_w*0 +:data_w] = c142obus[data_w*2 +:data_w];
assign c142ibus[temp_w*3 +:temp_w] = v727obus[temp_w*0 +:temp_w];
assign v727ibus[data_w*0 +:data_w] = c142obus[data_w*3 +:data_w];
assign c142ibus[temp_w*4 +:temp_w] = v1114obus[temp_w*0 +:temp_w];
assign v1114ibus[data_w*0 +:data_w] = c142obus[data_w*4 +:data_w];
assign c142ibus[temp_w*5 +:temp_w] = v1294obus[temp_w*1 +:temp_w];
assign v1294ibus[data_w*1 +:data_w] = c142obus[data_w*5 +:data_w];
assign c142ibus[temp_w*6 +:temp_w] = v1390obus[temp_w*0 +:temp_w];
assign v1390ibus[data_w*0 +:data_w] = c142obus[data_w*6 +:data_w];
assign c143ibus[temp_w*0 +:temp_w] = v170obus[temp_w*1 +:temp_w];
assign v170ibus[data_w*1 +:data_w] = c143obus[data_w*0 +:data_w];
assign c143ibus[temp_w*1 +:temp_w] = v549obus[temp_w*0 +:temp_w];
assign v549ibus[data_w*0 +:data_w] = c143obus[data_w*1 +:data_w];
assign c143ibus[temp_w*2 +:temp_w] = v606obus[temp_w*0 +:temp_w];
assign v606ibus[data_w*0 +:data_w] = c143obus[data_w*2 +:data_w];
assign c143ibus[temp_w*3 +:temp_w] = v728obus[temp_w*0 +:temp_w];
assign v728ibus[data_w*0 +:data_w] = c143obus[data_w*3 +:data_w];
assign c143ibus[temp_w*4 +:temp_w] = v1115obus[temp_w*0 +:temp_w];
assign v1115ibus[data_w*0 +:data_w] = c143obus[data_w*4 +:data_w];
assign c143ibus[temp_w*5 +:temp_w] = v1295obus[temp_w*1 +:temp_w];
assign v1295ibus[data_w*1 +:data_w] = c143obus[data_w*5 +:data_w];
assign c143ibus[temp_w*6 +:temp_w] = v1391obus[temp_w*0 +:temp_w];
assign v1391ibus[data_w*0 +:data_w] = c143obus[data_w*6 +:data_w];
assign c144ibus[temp_w*0 +:temp_w] = v171obus[temp_w*1 +:temp_w];
assign v171ibus[data_w*1 +:data_w] = c144obus[data_w*0 +:data_w];
assign c144ibus[temp_w*1 +:temp_w] = v550obus[temp_w*0 +:temp_w];
assign v550ibus[data_w*0 +:data_w] = c144obus[data_w*1 +:data_w];
assign c144ibus[temp_w*2 +:temp_w] = v607obus[temp_w*0 +:temp_w];
assign v607ibus[data_w*0 +:data_w] = c144obus[data_w*2 +:data_w];
assign c144ibus[temp_w*3 +:temp_w] = v729obus[temp_w*0 +:temp_w];
assign v729ibus[data_w*0 +:data_w] = c144obus[data_w*3 +:data_w];
assign c144ibus[temp_w*4 +:temp_w] = v1116obus[temp_w*0 +:temp_w];
assign v1116ibus[data_w*0 +:data_w] = c144obus[data_w*4 +:data_w];
assign c144ibus[temp_w*5 +:temp_w] = v1296obus[temp_w*1 +:temp_w];
assign v1296ibus[data_w*1 +:data_w] = c144obus[data_w*5 +:data_w];
assign c144ibus[temp_w*6 +:temp_w] = v1392obus[temp_w*0 +:temp_w];
assign v1392ibus[data_w*0 +:data_w] = c144obus[data_w*6 +:data_w];
assign c145ibus[temp_w*0 +:temp_w] = v172obus[temp_w*1 +:temp_w];
assign v172ibus[data_w*1 +:data_w] = c145obus[data_w*0 +:data_w];
assign c145ibus[temp_w*1 +:temp_w] = v551obus[temp_w*0 +:temp_w];
assign v551ibus[data_w*0 +:data_w] = c145obus[data_w*1 +:data_w];
assign c145ibus[temp_w*2 +:temp_w] = v608obus[temp_w*0 +:temp_w];
assign v608ibus[data_w*0 +:data_w] = c145obus[data_w*2 +:data_w];
assign c145ibus[temp_w*3 +:temp_w] = v730obus[temp_w*0 +:temp_w];
assign v730ibus[data_w*0 +:data_w] = c145obus[data_w*3 +:data_w];
assign c145ibus[temp_w*4 +:temp_w] = v1117obus[temp_w*0 +:temp_w];
assign v1117ibus[data_w*0 +:data_w] = c145obus[data_w*4 +:data_w];
assign c145ibus[temp_w*5 +:temp_w] = v1297obus[temp_w*1 +:temp_w];
assign v1297ibus[data_w*1 +:data_w] = c145obus[data_w*5 +:data_w];
assign c145ibus[temp_w*6 +:temp_w] = v1393obus[temp_w*0 +:temp_w];
assign v1393ibus[data_w*0 +:data_w] = c145obus[data_w*6 +:data_w];
assign c146ibus[temp_w*0 +:temp_w] = v173obus[temp_w*1 +:temp_w];
assign v173ibus[data_w*1 +:data_w] = c146obus[data_w*0 +:data_w];
assign c146ibus[temp_w*1 +:temp_w] = v552obus[temp_w*0 +:temp_w];
assign v552ibus[data_w*0 +:data_w] = c146obus[data_w*1 +:data_w];
assign c146ibus[temp_w*2 +:temp_w] = v609obus[temp_w*0 +:temp_w];
assign v609ibus[data_w*0 +:data_w] = c146obus[data_w*2 +:data_w];
assign c146ibus[temp_w*3 +:temp_w] = v731obus[temp_w*0 +:temp_w];
assign v731ibus[data_w*0 +:data_w] = c146obus[data_w*3 +:data_w];
assign c146ibus[temp_w*4 +:temp_w] = v1118obus[temp_w*0 +:temp_w];
assign v1118ibus[data_w*0 +:data_w] = c146obus[data_w*4 +:data_w];
assign c146ibus[temp_w*5 +:temp_w] = v1298obus[temp_w*1 +:temp_w];
assign v1298ibus[data_w*1 +:data_w] = c146obus[data_w*5 +:data_w];
assign c146ibus[temp_w*6 +:temp_w] = v1394obus[temp_w*0 +:temp_w];
assign v1394ibus[data_w*0 +:data_w] = c146obus[data_w*6 +:data_w];
assign c147ibus[temp_w*0 +:temp_w] = v174obus[temp_w*1 +:temp_w];
assign v174ibus[data_w*1 +:data_w] = c147obus[data_w*0 +:data_w];
assign c147ibus[temp_w*1 +:temp_w] = v553obus[temp_w*0 +:temp_w];
assign v553ibus[data_w*0 +:data_w] = c147obus[data_w*1 +:data_w];
assign c147ibus[temp_w*2 +:temp_w] = v610obus[temp_w*0 +:temp_w];
assign v610ibus[data_w*0 +:data_w] = c147obus[data_w*2 +:data_w];
assign c147ibus[temp_w*3 +:temp_w] = v732obus[temp_w*0 +:temp_w];
assign v732ibus[data_w*0 +:data_w] = c147obus[data_w*3 +:data_w];
assign c147ibus[temp_w*4 +:temp_w] = v1119obus[temp_w*0 +:temp_w];
assign v1119ibus[data_w*0 +:data_w] = c147obus[data_w*4 +:data_w];
assign c147ibus[temp_w*5 +:temp_w] = v1299obus[temp_w*1 +:temp_w];
assign v1299ibus[data_w*1 +:data_w] = c147obus[data_w*5 +:data_w];
assign c147ibus[temp_w*6 +:temp_w] = v1395obus[temp_w*0 +:temp_w];
assign v1395ibus[data_w*0 +:data_w] = c147obus[data_w*6 +:data_w];
assign c148ibus[temp_w*0 +:temp_w] = v175obus[temp_w*1 +:temp_w];
assign v175ibus[data_w*1 +:data_w] = c148obus[data_w*0 +:data_w];
assign c148ibus[temp_w*1 +:temp_w] = v554obus[temp_w*0 +:temp_w];
assign v554ibus[data_w*0 +:data_w] = c148obus[data_w*1 +:data_w];
assign c148ibus[temp_w*2 +:temp_w] = v611obus[temp_w*0 +:temp_w];
assign v611ibus[data_w*0 +:data_w] = c148obus[data_w*2 +:data_w];
assign c148ibus[temp_w*3 +:temp_w] = v733obus[temp_w*0 +:temp_w];
assign v733ibus[data_w*0 +:data_w] = c148obus[data_w*3 +:data_w];
assign c148ibus[temp_w*4 +:temp_w] = v1120obus[temp_w*0 +:temp_w];
assign v1120ibus[data_w*0 +:data_w] = c148obus[data_w*4 +:data_w];
assign c148ibus[temp_w*5 +:temp_w] = v1300obus[temp_w*1 +:temp_w];
assign v1300ibus[data_w*1 +:data_w] = c148obus[data_w*5 +:data_w];
assign c148ibus[temp_w*6 +:temp_w] = v1396obus[temp_w*0 +:temp_w];
assign v1396ibus[data_w*0 +:data_w] = c148obus[data_w*6 +:data_w];
assign c149ibus[temp_w*0 +:temp_w] = v176obus[temp_w*1 +:temp_w];
assign v176ibus[data_w*1 +:data_w] = c149obus[data_w*0 +:data_w];
assign c149ibus[temp_w*1 +:temp_w] = v555obus[temp_w*0 +:temp_w];
assign v555ibus[data_w*0 +:data_w] = c149obus[data_w*1 +:data_w];
assign c149ibus[temp_w*2 +:temp_w] = v612obus[temp_w*0 +:temp_w];
assign v612ibus[data_w*0 +:data_w] = c149obus[data_w*2 +:data_w];
assign c149ibus[temp_w*3 +:temp_w] = v734obus[temp_w*0 +:temp_w];
assign v734ibus[data_w*0 +:data_w] = c149obus[data_w*3 +:data_w];
assign c149ibus[temp_w*4 +:temp_w] = v1121obus[temp_w*0 +:temp_w];
assign v1121ibus[data_w*0 +:data_w] = c149obus[data_w*4 +:data_w];
assign c149ibus[temp_w*5 +:temp_w] = v1301obus[temp_w*1 +:temp_w];
assign v1301ibus[data_w*1 +:data_w] = c149obus[data_w*5 +:data_w];
assign c149ibus[temp_w*6 +:temp_w] = v1397obus[temp_w*0 +:temp_w];
assign v1397ibus[data_w*0 +:data_w] = c149obus[data_w*6 +:data_w];
assign c150ibus[temp_w*0 +:temp_w] = v177obus[temp_w*1 +:temp_w];
assign v177ibus[data_w*1 +:data_w] = c150obus[data_w*0 +:data_w];
assign c150ibus[temp_w*1 +:temp_w] = v556obus[temp_w*0 +:temp_w];
assign v556ibus[data_w*0 +:data_w] = c150obus[data_w*1 +:data_w];
assign c150ibus[temp_w*2 +:temp_w] = v613obus[temp_w*0 +:temp_w];
assign v613ibus[data_w*0 +:data_w] = c150obus[data_w*2 +:data_w];
assign c150ibus[temp_w*3 +:temp_w] = v735obus[temp_w*0 +:temp_w];
assign v735ibus[data_w*0 +:data_w] = c150obus[data_w*3 +:data_w];
assign c150ibus[temp_w*4 +:temp_w] = v1122obus[temp_w*0 +:temp_w];
assign v1122ibus[data_w*0 +:data_w] = c150obus[data_w*4 +:data_w];
assign c150ibus[temp_w*5 +:temp_w] = v1302obus[temp_w*1 +:temp_w];
assign v1302ibus[data_w*1 +:data_w] = c150obus[data_w*5 +:data_w];
assign c150ibus[temp_w*6 +:temp_w] = v1398obus[temp_w*0 +:temp_w];
assign v1398ibus[data_w*0 +:data_w] = c150obus[data_w*6 +:data_w];
assign c151ibus[temp_w*0 +:temp_w] = v178obus[temp_w*1 +:temp_w];
assign v178ibus[data_w*1 +:data_w] = c151obus[data_w*0 +:data_w];
assign c151ibus[temp_w*1 +:temp_w] = v557obus[temp_w*0 +:temp_w];
assign v557ibus[data_w*0 +:data_w] = c151obus[data_w*1 +:data_w];
assign c151ibus[temp_w*2 +:temp_w] = v614obus[temp_w*0 +:temp_w];
assign v614ibus[data_w*0 +:data_w] = c151obus[data_w*2 +:data_w];
assign c151ibus[temp_w*3 +:temp_w] = v736obus[temp_w*0 +:temp_w];
assign v736ibus[data_w*0 +:data_w] = c151obus[data_w*3 +:data_w];
assign c151ibus[temp_w*4 +:temp_w] = v1123obus[temp_w*0 +:temp_w];
assign v1123ibus[data_w*0 +:data_w] = c151obus[data_w*4 +:data_w];
assign c151ibus[temp_w*5 +:temp_w] = v1303obus[temp_w*1 +:temp_w];
assign v1303ibus[data_w*1 +:data_w] = c151obus[data_w*5 +:data_w];
assign c151ibus[temp_w*6 +:temp_w] = v1399obus[temp_w*0 +:temp_w];
assign v1399ibus[data_w*0 +:data_w] = c151obus[data_w*6 +:data_w];
assign c152ibus[temp_w*0 +:temp_w] = v179obus[temp_w*1 +:temp_w];
assign v179ibus[data_w*1 +:data_w] = c152obus[data_w*0 +:data_w];
assign c152ibus[temp_w*1 +:temp_w] = v558obus[temp_w*0 +:temp_w];
assign v558ibus[data_w*0 +:data_w] = c152obus[data_w*1 +:data_w];
assign c152ibus[temp_w*2 +:temp_w] = v615obus[temp_w*0 +:temp_w];
assign v615ibus[data_w*0 +:data_w] = c152obus[data_w*2 +:data_w];
assign c152ibus[temp_w*3 +:temp_w] = v737obus[temp_w*0 +:temp_w];
assign v737ibus[data_w*0 +:data_w] = c152obus[data_w*3 +:data_w];
assign c152ibus[temp_w*4 +:temp_w] = v1124obus[temp_w*0 +:temp_w];
assign v1124ibus[data_w*0 +:data_w] = c152obus[data_w*4 +:data_w];
assign c152ibus[temp_w*5 +:temp_w] = v1304obus[temp_w*1 +:temp_w];
assign v1304ibus[data_w*1 +:data_w] = c152obus[data_w*5 +:data_w];
assign c152ibus[temp_w*6 +:temp_w] = v1400obus[temp_w*0 +:temp_w];
assign v1400ibus[data_w*0 +:data_w] = c152obus[data_w*6 +:data_w];
assign c153ibus[temp_w*0 +:temp_w] = v180obus[temp_w*1 +:temp_w];
assign v180ibus[data_w*1 +:data_w] = c153obus[data_w*0 +:data_w];
assign c153ibus[temp_w*1 +:temp_w] = v559obus[temp_w*0 +:temp_w];
assign v559ibus[data_w*0 +:data_w] = c153obus[data_w*1 +:data_w];
assign c153ibus[temp_w*2 +:temp_w] = v616obus[temp_w*0 +:temp_w];
assign v616ibus[data_w*0 +:data_w] = c153obus[data_w*2 +:data_w];
assign c153ibus[temp_w*3 +:temp_w] = v738obus[temp_w*0 +:temp_w];
assign v738ibus[data_w*0 +:data_w] = c153obus[data_w*3 +:data_w];
assign c153ibus[temp_w*4 +:temp_w] = v1125obus[temp_w*0 +:temp_w];
assign v1125ibus[data_w*0 +:data_w] = c153obus[data_w*4 +:data_w];
assign c153ibus[temp_w*5 +:temp_w] = v1305obus[temp_w*1 +:temp_w];
assign v1305ibus[data_w*1 +:data_w] = c153obus[data_w*5 +:data_w];
assign c153ibus[temp_w*6 +:temp_w] = v1401obus[temp_w*0 +:temp_w];
assign v1401ibus[data_w*0 +:data_w] = c153obus[data_w*6 +:data_w];
assign c154ibus[temp_w*0 +:temp_w] = v181obus[temp_w*1 +:temp_w];
assign v181ibus[data_w*1 +:data_w] = c154obus[data_w*0 +:data_w];
assign c154ibus[temp_w*1 +:temp_w] = v560obus[temp_w*0 +:temp_w];
assign v560ibus[data_w*0 +:data_w] = c154obus[data_w*1 +:data_w];
assign c154ibus[temp_w*2 +:temp_w] = v617obus[temp_w*0 +:temp_w];
assign v617ibus[data_w*0 +:data_w] = c154obus[data_w*2 +:data_w];
assign c154ibus[temp_w*3 +:temp_w] = v739obus[temp_w*0 +:temp_w];
assign v739ibus[data_w*0 +:data_w] = c154obus[data_w*3 +:data_w];
assign c154ibus[temp_w*4 +:temp_w] = v1126obus[temp_w*0 +:temp_w];
assign v1126ibus[data_w*0 +:data_w] = c154obus[data_w*4 +:data_w];
assign c154ibus[temp_w*5 +:temp_w] = v1306obus[temp_w*1 +:temp_w];
assign v1306ibus[data_w*1 +:data_w] = c154obus[data_w*5 +:data_w];
assign c154ibus[temp_w*6 +:temp_w] = v1402obus[temp_w*0 +:temp_w];
assign v1402ibus[data_w*0 +:data_w] = c154obus[data_w*6 +:data_w];
assign c155ibus[temp_w*0 +:temp_w] = v182obus[temp_w*1 +:temp_w];
assign v182ibus[data_w*1 +:data_w] = c155obus[data_w*0 +:data_w];
assign c155ibus[temp_w*1 +:temp_w] = v561obus[temp_w*0 +:temp_w];
assign v561ibus[data_w*0 +:data_w] = c155obus[data_w*1 +:data_w];
assign c155ibus[temp_w*2 +:temp_w] = v618obus[temp_w*0 +:temp_w];
assign v618ibus[data_w*0 +:data_w] = c155obus[data_w*2 +:data_w];
assign c155ibus[temp_w*3 +:temp_w] = v740obus[temp_w*0 +:temp_w];
assign v740ibus[data_w*0 +:data_w] = c155obus[data_w*3 +:data_w];
assign c155ibus[temp_w*4 +:temp_w] = v1127obus[temp_w*0 +:temp_w];
assign v1127ibus[data_w*0 +:data_w] = c155obus[data_w*4 +:data_w];
assign c155ibus[temp_w*5 +:temp_w] = v1307obus[temp_w*1 +:temp_w];
assign v1307ibus[data_w*1 +:data_w] = c155obus[data_w*5 +:data_w];
assign c155ibus[temp_w*6 +:temp_w] = v1403obus[temp_w*0 +:temp_w];
assign v1403ibus[data_w*0 +:data_w] = c155obus[data_w*6 +:data_w];
assign c156ibus[temp_w*0 +:temp_w] = v183obus[temp_w*1 +:temp_w];
assign v183ibus[data_w*1 +:data_w] = c156obus[data_w*0 +:data_w];
assign c156ibus[temp_w*1 +:temp_w] = v562obus[temp_w*0 +:temp_w];
assign v562ibus[data_w*0 +:data_w] = c156obus[data_w*1 +:data_w];
assign c156ibus[temp_w*2 +:temp_w] = v619obus[temp_w*0 +:temp_w];
assign v619ibus[data_w*0 +:data_w] = c156obus[data_w*2 +:data_w];
assign c156ibus[temp_w*3 +:temp_w] = v741obus[temp_w*0 +:temp_w];
assign v741ibus[data_w*0 +:data_w] = c156obus[data_w*3 +:data_w];
assign c156ibus[temp_w*4 +:temp_w] = v1128obus[temp_w*0 +:temp_w];
assign v1128ibus[data_w*0 +:data_w] = c156obus[data_w*4 +:data_w];
assign c156ibus[temp_w*5 +:temp_w] = v1308obus[temp_w*1 +:temp_w];
assign v1308ibus[data_w*1 +:data_w] = c156obus[data_w*5 +:data_w];
assign c156ibus[temp_w*6 +:temp_w] = v1404obus[temp_w*0 +:temp_w];
assign v1404ibus[data_w*0 +:data_w] = c156obus[data_w*6 +:data_w];
assign c157ibus[temp_w*0 +:temp_w] = v184obus[temp_w*1 +:temp_w];
assign v184ibus[data_w*1 +:data_w] = c157obus[data_w*0 +:data_w];
assign c157ibus[temp_w*1 +:temp_w] = v563obus[temp_w*0 +:temp_w];
assign v563ibus[data_w*0 +:data_w] = c157obus[data_w*1 +:data_w];
assign c157ibus[temp_w*2 +:temp_w] = v620obus[temp_w*0 +:temp_w];
assign v620ibus[data_w*0 +:data_w] = c157obus[data_w*2 +:data_w];
assign c157ibus[temp_w*3 +:temp_w] = v742obus[temp_w*0 +:temp_w];
assign v742ibus[data_w*0 +:data_w] = c157obus[data_w*3 +:data_w];
assign c157ibus[temp_w*4 +:temp_w] = v1129obus[temp_w*0 +:temp_w];
assign v1129ibus[data_w*0 +:data_w] = c157obus[data_w*4 +:data_w];
assign c157ibus[temp_w*5 +:temp_w] = v1309obus[temp_w*1 +:temp_w];
assign v1309ibus[data_w*1 +:data_w] = c157obus[data_w*5 +:data_w];
assign c157ibus[temp_w*6 +:temp_w] = v1405obus[temp_w*0 +:temp_w];
assign v1405ibus[data_w*0 +:data_w] = c157obus[data_w*6 +:data_w];
assign c158ibus[temp_w*0 +:temp_w] = v185obus[temp_w*1 +:temp_w];
assign v185ibus[data_w*1 +:data_w] = c158obus[data_w*0 +:data_w];
assign c158ibus[temp_w*1 +:temp_w] = v564obus[temp_w*0 +:temp_w];
assign v564ibus[data_w*0 +:data_w] = c158obus[data_w*1 +:data_w];
assign c158ibus[temp_w*2 +:temp_w] = v621obus[temp_w*0 +:temp_w];
assign v621ibus[data_w*0 +:data_w] = c158obus[data_w*2 +:data_w];
assign c158ibus[temp_w*3 +:temp_w] = v743obus[temp_w*0 +:temp_w];
assign v743ibus[data_w*0 +:data_w] = c158obus[data_w*3 +:data_w];
assign c158ibus[temp_w*4 +:temp_w] = v1130obus[temp_w*0 +:temp_w];
assign v1130ibus[data_w*0 +:data_w] = c158obus[data_w*4 +:data_w];
assign c158ibus[temp_w*5 +:temp_w] = v1310obus[temp_w*1 +:temp_w];
assign v1310ibus[data_w*1 +:data_w] = c158obus[data_w*5 +:data_w];
assign c158ibus[temp_w*6 +:temp_w] = v1406obus[temp_w*0 +:temp_w];
assign v1406ibus[data_w*0 +:data_w] = c158obus[data_w*6 +:data_w];
assign c159ibus[temp_w*0 +:temp_w] = v186obus[temp_w*1 +:temp_w];
assign v186ibus[data_w*1 +:data_w] = c159obus[data_w*0 +:data_w];
assign c159ibus[temp_w*1 +:temp_w] = v565obus[temp_w*0 +:temp_w];
assign v565ibus[data_w*0 +:data_w] = c159obus[data_w*1 +:data_w];
assign c159ibus[temp_w*2 +:temp_w] = v622obus[temp_w*0 +:temp_w];
assign v622ibus[data_w*0 +:data_w] = c159obus[data_w*2 +:data_w];
assign c159ibus[temp_w*3 +:temp_w] = v744obus[temp_w*0 +:temp_w];
assign v744ibus[data_w*0 +:data_w] = c159obus[data_w*3 +:data_w];
assign c159ibus[temp_w*4 +:temp_w] = v1131obus[temp_w*0 +:temp_w];
assign v1131ibus[data_w*0 +:data_w] = c159obus[data_w*4 +:data_w];
assign c159ibus[temp_w*5 +:temp_w] = v1311obus[temp_w*1 +:temp_w];
assign v1311ibus[data_w*1 +:data_w] = c159obus[data_w*5 +:data_w];
assign c159ibus[temp_w*6 +:temp_w] = v1407obus[temp_w*0 +:temp_w];
assign v1407ibus[data_w*0 +:data_w] = c159obus[data_w*6 +:data_w];
assign c160ibus[temp_w*0 +:temp_w] = v187obus[temp_w*1 +:temp_w];
assign v187ibus[data_w*1 +:data_w] = c160obus[data_w*0 +:data_w];
assign c160ibus[temp_w*1 +:temp_w] = v566obus[temp_w*0 +:temp_w];
assign v566ibus[data_w*0 +:data_w] = c160obus[data_w*1 +:data_w];
assign c160ibus[temp_w*2 +:temp_w] = v623obus[temp_w*0 +:temp_w];
assign v623ibus[data_w*0 +:data_w] = c160obus[data_w*2 +:data_w];
assign c160ibus[temp_w*3 +:temp_w] = v745obus[temp_w*0 +:temp_w];
assign v745ibus[data_w*0 +:data_w] = c160obus[data_w*3 +:data_w];
assign c160ibus[temp_w*4 +:temp_w] = v1132obus[temp_w*0 +:temp_w];
assign v1132ibus[data_w*0 +:data_w] = c160obus[data_w*4 +:data_w];
assign c160ibus[temp_w*5 +:temp_w] = v1312obus[temp_w*1 +:temp_w];
assign v1312ibus[data_w*1 +:data_w] = c160obus[data_w*5 +:data_w];
assign c160ibus[temp_w*6 +:temp_w] = v1408obus[temp_w*0 +:temp_w];
assign v1408ibus[data_w*0 +:data_w] = c160obus[data_w*6 +:data_w];
assign c161ibus[temp_w*0 +:temp_w] = v188obus[temp_w*1 +:temp_w];
assign v188ibus[data_w*1 +:data_w] = c161obus[data_w*0 +:data_w];
assign c161ibus[temp_w*1 +:temp_w] = v567obus[temp_w*0 +:temp_w];
assign v567ibus[data_w*0 +:data_w] = c161obus[data_w*1 +:data_w];
assign c161ibus[temp_w*2 +:temp_w] = v624obus[temp_w*0 +:temp_w];
assign v624ibus[data_w*0 +:data_w] = c161obus[data_w*2 +:data_w];
assign c161ibus[temp_w*3 +:temp_w] = v746obus[temp_w*0 +:temp_w];
assign v746ibus[data_w*0 +:data_w] = c161obus[data_w*3 +:data_w];
assign c161ibus[temp_w*4 +:temp_w] = v1133obus[temp_w*0 +:temp_w];
assign v1133ibus[data_w*0 +:data_w] = c161obus[data_w*4 +:data_w];
assign c161ibus[temp_w*5 +:temp_w] = v1313obus[temp_w*1 +:temp_w];
assign v1313ibus[data_w*1 +:data_w] = c161obus[data_w*5 +:data_w];
assign c161ibus[temp_w*6 +:temp_w] = v1409obus[temp_w*0 +:temp_w];
assign v1409ibus[data_w*0 +:data_w] = c161obus[data_w*6 +:data_w];
assign c162ibus[temp_w*0 +:temp_w] = v189obus[temp_w*1 +:temp_w];
assign v189ibus[data_w*1 +:data_w] = c162obus[data_w*0 +:data_w];
assign c162ibus[temp_w*1 +:temp_w] = v568obus[temp_w*0 +:temp_w];
assign v568ibus[data_w*0 +:data_w] = c162obus[data_w*1 +:data_w];
assign c162ibus[temp_w*2 +:temp_w] = v625obus[temp_w*0 +:temp_w];
assign v625ibus[data_w*0 +:data_w] = c162obus[data_w*2 +:data_w];
assign c162ibus[temp_w*3 +:temp_w] = v747obus[temp_w*0 +:temp_w];
assign v747ibus[data_w*0 +:data_w] = c162obus[data_w*3 +:data_w];
assign c162ibus[temp_w*4 +:temp_w] = v1134obus[temp_w*0 +:temp_w];
assign v1134ibus[data_w*0 +:data_w] = c162obus[data_w*4 +:data_w];
assign c162ibus[temp_w*5 +:temp_w] = v1314obus[temp_w*1 +:temp_w];
assign v1314ibus[data_w*1 +:data_w] = c162obus[data_w*5 +:data_w];
assign c162ibus[temp_w*6 +:temp_w] = v1410obus[temp_w*0 +:temp_w];
assign v1410ibus[data_w*0 +:data_w] = c162obus[data_w*6 +:data_w];
assign c163ibus[temp_w*0 +:temp_w] = v190obus[temp_w*1 +:temp_w];
assign v190ibus[data_w*1 +:data_w] = c163obus[data_w*0 +:data_w];
assign c163ibus[temp_w*1 +:temp_w] = v569obus[temp_w*0 +:temp_w];
assign v569ibus[data_w*0 +:data_w] = c163obus[data_w*1 +:data_w];
assign c163ibus[temp_w*2 +:temp_w] = v626obus[temp_w*0 +:temp_w];
assign v626ibus[data_w*0 +:data_w] = c163obus[data_w*2 +:data_w];
assign c163ibus[temp_w*3 +:temp_w] = v748obus[temp_w*0 +:temp_w];
assign v748ibus[data_w*0 +:data_w] = c163obus[data_w*3 +:data_w];
assign c163ibus[temp_w*4 +:temp_w] = v1135obus[temp_w*0 +:temp_w];
assign v1135ibus[data_w*0 +:data_w] = c163obus[data_w*4 +:data_w];
assign c163ibus[temp_w*5 +:temp_w] = v1315obus[temp_w*1 +:temp_w];
assign v1315ibus[data_w*1 +:data_w] = c163obus[data_w*5 +:data_w];
assign c163ibus[temp_w*6 +:temp_w] = v1411obus[temp_w*0 +:temp_w];
assign v1411ibus[data_w*0 +:data_w] = c163obus[data_w*6 +:data_w];
assign c164ibus[temp_w*0 +:temp_w] = v191obus[temp_w*1 +:temp_w];
assign v191ibus[data_w*1 +:data_w] = c164obus[data_w*0 +:data_w];
assign c164ibus[temp_w*1 +:temp_w] = v570obus[temp_w*0 +:temp_w];
assign v570ibus[data_w*0 +:data_w] = c164obus[data_w*1 +:data_w];
assign c164ibus[temp_w*2 +:temp_w] = v627obus[temp_w*0 +:temp_w];
assign v627ibus[data_w*0 +:data_w] = c164obus[data_w*2 +:data_w];
assign c164ibus[temp_w*3 +:temp_w] = v749obus[temp_w*0 +:temp_w];
assign v749ibus[data_w*0 +:data_w] = c164obus[data_w*3 +:data_w];
assign c164ibus[temp_w*4 +:temp_w] = v1136obus[temp_w*0 +:temp_w];
assign v1136ibus[data_w*0 +:data_w] = c164obus[data_w*4 +:data_w];
assign c164ibus[temp_w*5 +:temp_w] = v1316obus[temp_w*1 +:temp_w];
assign v1316ibus[data_w*1 +:data_w] = c164obus[data_w*5 +:data_w];
assign c164ibus[temp_w*6 +:temp_w] = v1412obus[temp_w*0 +:temp_w];
assign v1412ibus[data_w*0 +:data_w] = c164obus[data_w*6 +:data_w];
assign c165ibus[temp_w*0 +:temp_w] = v96obus[temp_w*1 +:temp_w];
assign v96ibus[data_w*1 +:data_w] = c165obus[data_w*0 +:data_w];
assign c165ibus[temp_w*1 +:temp_w] = v571obus[temp_w*0 +:temp_w];
assign v571ibus[data_w*0 +:data_w] = c165obus[data_w*1 +:data_w];
assign c165ibus[temp_w*2 +:temp_w] = v628obus[temp_w*0 +:temp_w];
assign v628ibus[data_w*0 +:data_w] = c165obus[data_w*2 +:data_w];
assign c165ibus[temp_w*3 +:temp_w] = v750obus[temp_w*0 +:temp_w];
assign v750ibus[data_w*0 +:data_w] = c165obus[data_w*3 +:data_w];
assign c165ibus[temp_w*4 +:temp_w] = v1137obus[temp_w*0 +:temp_w];
assign v1137ibus[data_w*0 +:data_w] = c165obus[data_w*4 +:data_w];
assign c165ibus[temp_w*5 +:temp_w] = v1317obus[temp_w*1 +:temp_w];
assign v1317ibus[data_w*1 +:data_w] = c165obus[data_w*5 +:data_w];
assign c165ibus[temp_w*6 +:temp_w] = v1413obus[temp_w*0 +:temp_w];
assign v1413ibus[data_w*0 +:data_w] = c165obus[data_w*6 +:data_w];
assign c166ibus[temp_w*0 +:temp_w] = v97obus[temp_w*1 +:temp_w];
assign v97ibus[data_w*1 +:data_w] = c166obus[data_w*0 +:data_w];
assign c166ibus[temp_w*1 +:temp_w] = v572obus[temp_w*0 +:temp_w];
assign v572ibus[data_w*0 +:data_w] = c166obus[data_w*1 +:data_w];
assign c166ibus[temp_w*2 +:temp_w] = v629obus[temp_w*0 +:temp_w];
assign v629ibus[data_w*0 +:data_w] = c166obus[data_w*2 +:data_w];
assign c166ibus[temp_w*3 +:temp_w] = v751obus[temp_w*0 +:temp_w];
assign v751ibus[data_w*0 +:data_w] = c166obus[data_w*3 +:data_w];
assign c166ibus[temp_w*4 +:temp_w] = v1138obus[temp_w*0 +:temp_w];
assign v1138ibus[data_w*0 +:data_w] = c166obus[data_w*4 +:data_w];
assign c166ibus[temp_w*5 +:temp_w] = v1318obus[temp_w*1 +:temp_w];
assign v1318ibus[data_w*1 +:data_w] = c166obus[data_w*5 +:data_w];
assign c166ibus[temp_w*6 +:temp_w] = v1414obus[temp_w*0 +:temp_w];
assign v1414ibus[data_w*0 +:data_w] = c166obus[data_w*6 +:data_w];
assign c167ibus[temp_w*0 +:temp_w] = v98obus[temp_w*1 +:temp_w];
assign v98ibus[data_w*1 +:data_w] = c167obus[data_w*0 +:data_w];
assign c167ibus[temp_w*1 +:temp_w] = v573obus[temp_w*0 +:temp_w];
assign v573ibus[data_w*0 +:data_w] = c167obus[data_w*1 +:data_w];
assign c167ibus[temp_w*2 +:temp_w] = v630obus[temp_w*0 +:temp_w];
assign v630ibus[data_w*0 +:data_w] = c167obus[data_w*2 +:data_w];
assign c167ibus[temp_w*3 +:temp_w] = v752obus[temp_w*0 +:temp_w];
assign v752ibus[data_w*0 +:data_w] = c167obus[data_w*3 +:data_w];
assign c167ibus[temp_w*4 +:temp_w] = v1139obus[temp_w*0 +:temp_w];
assign v1139ibus[data_w*0 +:data_w] = c167obus[data_w*4 +:data_w];
assign c167ibus[temp_w*5 +:temp_w] = v1319obus[temp_w*1 +:temp_w];
assign v1319ibus[data_w*1 +:data_w] = c167obus[data_w*5 +:data_w];
assign c167ibus[temp_w*6 +:temp_w] = v1415obus[temp_w*0 +:temp_w];
assign v1415ibus[data_w*0 +:data_w] = c167obus[data_w*6 +:data_w];
assign c168ibus[temp_w*0 +:temp_w] = v99obus[temp_w*1 +:temp_w];
assign v99ibus[data_w*1 +:data_w] = c168obus[data_w*0 +:data_w];
assign c168ibus[temp_w*1 +:temp_w] = v574obus[temp_w*0 +:temp_w];
assign v574ibus[data_w*0 +:data_w] = c168obus[data_w*1 +:data_w];
assign c168ibus[temp_w*2 +:temp_w] = v631obus[temp_w*0 +:temp_w];
assign v631ibus[data_w*0 +:data_w] = c168obus[data_w*2 +:data_w];
assign c168ibus[temp_w*3 +:temp_w] = v753obus[temp_w*0 +:temp_w];
assign v753ibus[data_w*0 +:data_w] = c168obus[data_w*3 +:data_w];
assign c168ibus[temp_w*4 +:temp_w] = v1140obus[temp_w*0 +:temp_w];
assign v1140ibus[data_w*0 +:data_w] = c168obus[data_w*4 +:data_w];
assign c168ibus[temp_w*5 +:temp_w] = v1320obus[temp_w*1 +:temp_w];
assign v1320ibus[data_w*1 +:data_w] = c168obus[data_w*5 +:data_w];
assign c168ibus[temp_w*6 +:temp_w] = v1416obus[temp_w*0 +:temp_w];
assign v1416ibus[data_w*0 +:data_w] = c168obus[data_w*6 +:data_w];
assign c169ibus[temp_w*0 +:temp_w] = v100obus[temp_w*1 +:temp_w];
assign v100ibus[data_w*1 +:data_w] = c169obus[data_w*0 +:data_w];
assign c169ibus[temp_w*1 +:temp_w] = v575obus[temp_w*0 +:temp_w];
assign v575ibus[data_w*0 +:data_w] = c169obus[data_w*1 +:data_w];
assign c169ibus[temp_w*2 +:temp_w] = v632obus[temp_w*0 +:temp_w];
assign v632ibus[data_w*0 +:data_w] = c169obus[data_w*2 +:data_w];
assign c169ibus[temp_w*3 +:temp_w] = v754obus[temp_w*0 +:temp_w];
assign v754ibus[data_w*0 +:data_w] = c169obus[data_w*3 +:data_w];
assign c169ibus[temp_w*4 +:temp_w] = v1141obus[temp_w*0 +:temp_w];
assign v1141ibus[data_w*0 +:data_w] = c169obus[data_w*4 +:data_w];
assign c169ibus[temp_w*5 +:temp_w] = v1321obus[temp_w*1 +:temp_w];
assign v1321ibus[data_w*1 +:data_w] = c169obus[data_w*5 +:data_w];
assign c169ibus[temp_w*6 +:temp_w] = v1417obus[temp_w*0 +:temp_w];
assign v1417ibus[data_w*0 +:data_w] = c169obus[data_w*6 +:data_w];
assign c170ibus[temp_w*0 +:temp_w] = v101obus[temp_w*1 +:temp_w];
assign v101ibus[data_w*1 +:data_w] = c170obus[data_w*0 +:data_w];
assign c170ibus[temp_w*1 +:temp_w] = v480obus[temp_w*0 +:temp_w];
assign v480ibus[data_w*0 +:data_w] = c170obus[data_w*1 +:data_w];
assign c170ibus[temp_w*2 +:temp_w] = v633obus[temp_w*0 +:temp_w];
assign v633ibus[data_w*0 +:data_w] = c170obus[data_w*2 +:data_w];
assign c170ibus[temp_w*3 +:temp_w] = v755obus[temp_w*0 +:temp_w];
assign v755ibus[data_w*0 +:data_w] = c170obus[data_w*3 +:data_w];
assign c170ibus[temp_w*4 +:temp_w] = v1142obus[temp_w*0 +:temp_w];
assign v1142ibus[data_w*0 +:data_w] = c170obus[data_w*4 +:data_w];
assign c170ibus[temp_w*5 +:temp_w] = v1322obus[temp_w*1 +:temp_w];
assign v1322ibus[data_w*1 +:data_w] = c170obus[data_w*5 +:data_w];
assign c170ibus[temp_w*6 +:temp_w] = v1418obus[temp_w*0 +:temp_w];
assign v1418ibus[data_w*0 +:data_w] = c170obus[data_w*6 +:data_w];
assign c171ibus[temp_w*0 +:temp_w] = v102obus[temp_w*1 +:temp_w];
assign v102ibus[data_w*1 +:data_w] = c171obus[data_w*0 +:data_w];
assign c171ibus[temp_w*1 +:temp_w] = v481obus[temp_w*0 +:temp_w];
assign v481ibus[data_w*0 +:data_w] = c171obus[data_w*1 +:data_w];
assign c171ibus[temp_w*2 +:temp_w] = v634obus[temp_w*0 +:temp_w];
assign v634ibus[data_w*0 +:data_w] = c171obus[data_w*2 +:data_w];
assign c171ibus[temp_w*3 +:temp_w] = v756obus[temp_w*0 +:temp_w];
assign v756ibus[data_w*0 +:data_w] = c171obus[data_w*3 +:data_w];
assign c171ibus[temp_w*4 +:temp_w] = v1143obus[temp_w*0 +:temp_w];
assign v1143ibus[data_w*0 +:data_w] = c171obus[data_w*4 +:data_w];
assign c171ibus[temp_w*5 +:temp_w] = v1323obus[temp_w*1 +:temp_w];
assign v1323ibus[data_w*1 +:data_w] = c171obus[data_w*5 +:data_w];
assign c171ibus[temp_w*6 +:temp_w] = v1419obus[temp_w*0 +:temp_w];
assign v1419ibus[data_w*0 +:data_w] = c171obus[data_w*6 +:data_w];
assign c172ibus[temp_w*0 +:temp_w] = v103obus[temp_w*1 +:temp_w];
assign v103ibus[data_w*1 +:data_w] = c172obus[data_w*0 +:data_w];
assign c172ibus[temp_w*1 +:temp_w] = v482obus[temp_w*0 +:temp_w];
assign v482ibus[data_w*0 +:data_w] = c172obus[data_w*1 +:data_w];
assign c172ibus[temp_w*2 +:temp_w] = v635obus[temp_w*0 +:temp_w];
assign v635ibus[data_w*0 +:data_w] = c172obus[data_w*2 +:data_w];
assign c172ibus[temp_w*3 +:temp_w] = v757obus[temp_w*0 +:temp_w];
assign v757ibus[data_w*0 +:data_w] = c172obus[data_w*3 +:data_w];
assign c172ibus[temp_w*4 +:temp_w] = v1144obus[temp_w*0 +:temp_w];
assign v1144ibus[data_w*0 +:data_w] = c172obus[data_w*4 +:data_w];
assign c172ibus[temp_w*5 +:temp_w] = v1324obus[temp_w*1 +:temp_w];
assign v1324ibus[data_w*1 +:data_w] = c172obus[data_w*5 +:data_w];
assign c172ibus[temp_w*6 +:temp_w] = v1420obus[temp_w*0 +:temp_w];
assign v1420ibus[data_w*0 +:data_w] = c172obus[data_w*6 +:data_w];
assign c173ibus[temp_w*0 +:temp_w] = v104obus[temp_w*1 +:temp_w];
assign v104ibus[data_w*1 +:data_w] = c173obus[data_w*0 +:data_w];
assign c173ibus[temp_w*1 +:temp_w] = v483obus[temp_w*0 +:temp_w];
assign v483ibus[data_w*0 +:data_w] = c173obus[data_w*1 +:data_w];
assign c173ibus[temp_w*2 +:temp_w] = v636obus[temp_w*0 +:temp_w];
assign v636ibus[data_w*0 +:data_w] = c173obus[data_w*2 +:data_w];
assign c173ibus[temp_w*3 +:temp_w] = v758obus[temp_w*0 +:temp_w];
assign v758ibus[data_w*0 +:data_w] = c173obus[data_w*3 +:data_w];
assign c173ibus[temp_w*4 +:temp_w] = v1145obus[temp_w*0 +:temp_w];
assign v1145ibus[data_w*0 +:data_w] = c173obus[data_w*4 +:data_w];
assign c173ibus[temp_w*5 +:temp_w] = v1325obus[temp_w*1 +:temp_w];
assign v1325ibus[data_w*1 +:data_w] = c173obus[data_w*5 +:data_w];
assign c173ibus[temp_w*6 +:temp_w] = v1421obus[temp_w*0 +:temp_w];
assign v1421ibus[data_w*0 +:data_w] = c173obus[data_w*6 +:data_w];
assign c174ibus[temp_w*0 +:temp_w] = v105obus[temp_w*1 +:temp_w];
assign v105ibus[data_w*1 +:data_w] = c174obus[data_w*0 +:data_w];
assign c174ibus[temp_w*1 +:temp_w] = v484obus[temp_w*0 +:temp_w];
assign v484ibus[data_w*0 +:data_w] = c174obus[data_w*1 +:data_w];
assign c174ibus[temp_w*2 +:temp_w] = v637obus[temp_w*0 +:temp_w];
assign v637ibus[data_w*0 +:data_w] = c174obus[data_w*2 +:data_w];
assign c174ibus[temp_w*3 +:temp_w] = v759obus[temp_w*0 +:temp_w];
assign v759ibus[data_w*0 +:data_w] = c174obus[data_w*3 +:data_w];
assign c174ibus[temp_w*4 +:temp_w] = v1146obus[temp_w*0 +:temp_w];
assign v1146ibus[data_w*0 +:data_w] = c174obus[data_w*4 +:data_w];
assign c174ibus[temp_w*5 +:temp_w] = v1326obus[temp_w*1 +:temp_w];
assign v1326ibus[data_w*1 +:data_w] = c174obus[data_w*5 +:data_w];
assign c174ibus[temp_w*6 +:temp_w] = v1422obus[temp_w*0 +:temp_w];
assign v1422ibus[data_w*0 +:data_w] = c174obus[data_w*6 +:data_w];
assign c175ibus[temp_w*0 +:temp_w] = v106obus[temp_w*1 +:temp_w];
assign v106ibus[data_w*1 +:data_w] = c175obus[data_w*0 +:data_w];
assign c175ibus[temp_w*1 +:temp_w] = v485obus[temp_w*0 +:temp_w];
assign v485ibus[data_w*0 +:data_w] = c175obus[data_w*1 +:data_w];
assign c175ibus[temp_w*2 +:temp_w] = v638obus[temp_w*0 +:temp_w];
assign v638ibus[data_w*0 +:data_w] = c175obus[data_w*2 +:data_w];
assign c175ibus[temp_w*3 +:temp_w] = v760obus[temp_w*0 +:temp_w];
assign v760ibus[data_w*0 +:data_w] = c175obus[data_w*3 +:data_w];
assign c175ibus[temp_w*4 +:temp_w] = v1147obus[temp_w*0 +:temp_w];
assign v1147ibus[data_w*0 +:data_w] = c175obus[data_w*4 +:data_w];
assign c175ibus[temp_w*5 +:temp_w] = v1327obus[temp_w*1 +:temp_w];
assign v1327ibus[data_w*1 +:data_w] = c175obus[data_w*5 +:data_w];
assign c175ibus[temp_w*6 +:temp_w] = v1423obus[temp_w*0 +:temp_w];
assign v1423ibus[data_w*0 +:data_w] = c175obus[data_w*6 +:data_w];
assign c176ibus[temp_w*0 +:temp_w] = v107obus[temp_w*1 +:temp_w];
assign v107ibus[data_w*1 +:data_w] = c176obus[data_w*0 +:data_w];
assign c176ibus[temp_w*1 +:temp_w] = v486obus[temp_w*0 +:temp_w];
assign v486ibus[data_w*0 +:data_w] = c176obus[data_w*1 +:data_w];
assign c176ibus[temp_w*2 +:temp_w] = v639obus[temp_w*0 +:temp_w];
assign v639ibus[data_w*0 +:data_w] = c176obus[data_w*2 +:data_w];
assign c176ibus[temp_w*3 +:temp_w] = v761obus[temp_w*0 +:temp_w];
assign v761ibus[data_w*0 +:data_w] = c176obus[data_w*3 +:data_w];
assign c176ibus[temp_w*4 +:temp_w] = v1148obus[temp_w*0 +:temp_w];
assign v1148ibus[data_w*0 +:data_w] = c176obus[data_w*4 +:data_w];
assign c176ibus[temp_w*5 +:temp_w] = v1328obus[temp_w*1 +:temp_w];
assign v1328ibus[data_w*1 +:data_w] = c176obus[data_w*5 +:data_w];
assign c176ibus[temp_w*6 +:temp_w] = v1424obus[temp_w*0 +:temp_w];
assign v1424ibus[data_w*0 +:data_w] = c176obus[data_w*6 +:data_w];
assign c177ibus[temp_w*0 +:temp_w] = v108obus[temp_w*1 +:temp_w];
assign v108ibus[data_w*1 +:data_w] = c177obus[data_w*0 +:data_w];
assign c177ibus[temp_w*1 +:temp_w] = v487obus[temp_w*0 +:temp_w];
assign v487ibus[data_w*0 +:data_w] = c177obus[data_w*1 +:data_w];
assign c177ibus[temp_w*2 +:temp_w] = v640obus[temp_w*0 +:temp_w];
assign v640ibus[data_w*0 +:data_w] = c177obus[data_w*2 +:data_w];
assign c177ibus[temp_w*3 +:temp_w] = v762obus[temp_w*0 +:temp_w];
assign v762ibus[data_w*0 +:data_w] = c177obus[data_w*3 +:data_w];
assign c177ibus[temp_w*4 +:temp_w] = v1149obus[temp_w*0 +:temp_w];
assign v1149ibus[data_w*0 +:data_w] = c177obus[data_w*4 +:data_w];
assign c177ibus[temp_w*5 +:temp_w] = v1329obus[temp_w*1 +:temp_w];
assign v1329ibus[data_w*1 +:data_w] = c177obus[data_w*5 +:data_w];
assign c177ibus[temp_w*6 +:temp_w] = v1425obus[temp_w*0 +:temp_w];
assign v1425ibus[data_w*0 +:data_w] = c177obus[data_w*6 +:data_w];
assign c178ibus[temp_w*0 +:temp_w] = v109obus[temp_w*1 +:temp_w];
assign v109ibus[data_w*1 +:data_w] = c178obus[data_w*0 +:data_w];
assign c178ibus[temp_w*1 +:temp_w] = v488obus[temp_w*0 +:temp_w];
assign v488ibus[data_w*0 +:data_w] = c178obus[data_w*1 +:data_w];
assign c178ibus[temp_w*2 +:temp_w] = v641obus[temp_w*0 +:temp_w];
assign v641ibus[data_w*0 +:data_w] = c178obus[data_w*2 +:data_w];
assign c178ibus[temp_w*3 +:temp_w] = v763obus[temp_w*0 +:temp_w];
assign v763ibus[data_w*0 +:data_w] = c178obus[data_w*3 +:data_w];
assign c178ibus[temp_w*4 +:temp_w] = v1150obus[temp_w*0 +:temp_w];
assign v1150ibus[data_w*0 +:data_w] = c178obus[data_w*4 +:data_w];
assign c178ibus[temp_w*5 +:temp_w] = v1330obus[temp_w*1 +:temp_w];
assign v1330ibus[data_w*1 +:data_w] = c178obus[data_w*5 +:data_w];
assign c178ibus[temp_w*6 +:temp_w] = v1426obus[temp_w*0 +:temp_w];
assign v1426ibus[data_w*0 +:data_w] = c178obus[data_w*6 +:data_w];
assign c179ibus[temp_w*0 +:temp_w] = v110obus[temp_w*1 +:temp_w];
assign v110ibus[data_w*1 +:data_w] = c179obus[data_w*0 +:data_w];
assign c179ibus[temp_w*1 +:temp_w] = v489obus[temp_w*0 +:temp_w];
assign v489ibus[data_w*0 +:data_w] = c179obus[data_w*1 +:data_w];
assign c179ibus[temp_w*2 +:temp_w] = v642obus[temp_w*0 +:temp_w];
assign v642ibus[data_w*0 +:data_w] = c179obus[data_w*2 +:data_w];
assign c179ibus[temp_w*3 +:temp_w] = v764obus[temp_w*0 +:temp_w];
assign v764ibus[data_w*0 +:data_w] = c179obus[data_w*3 +:data_w];
assign c179ibus[temp_w*4 +:temp_w] = v1151obus[temp_w*0 +:temp_w];
assign v1151ibus[data_w*0 +:data_w] = c179obus[data_w*4 +:data_w];
assign c179ibus[temp_w*5 +:temp_w] = v1331obus[temp_w*1 +:temp_w];
assign v1331ibus[data_w*1 +:data_w] = c179obus[data_w*5 +:data_w];
assign c179ibus[temp_w*6 +:temp_w] = v1427obus[temp_w*0 +:temp_w];
assign v1427ibus[data_w*0 +:data_w] = c179obus[data_w*6 +:data_w];
assign c180ibus[temp_w*0 +:temp_w] = v111obus[temp_w*1 +:temp_w];
assign v111ibus[data_w*1 +:data_w] = c180obus[data_w*0 +:data_w];
assign c180ibus[temp_w*1 +:temp_w] = v490obus[temp_w*0 +:temp_w];
assign v490ibus[data_w*0 +:data_w] = c180obus[data_w*1 +:data_w];
assign c180ibus[temp_w*2 +:temp_w] = v643obus[temp_w*0 +:temp_w];
assign v643ibus[data_w*0 +:data_w] = c180obus[data_w*2 +:data_w];
assign c180ibus[temp_w*3 +:temp_w] = v765obus[temp_w*0 +:temp_w];
assign v765ibus[data_w*0 +:data_w] = c180obus[data_w*3 +:data_w];
assign c180ibus[temp_w*4 +:temp_w] = v1056obus[temp_w*0 +:temp_w];
assign v1056ibus[data_w*0 +:data_w] = c180obus[data_w*4 +:data_w];
assign c180ibus[temp_w*5 +:temp_w] = v1332obus[temp_w*1 +:temp_w];
assign v1332ibus[data_w*1 +:data_w] = c180obus[data_w*5 +:data_w];
assign c180ibus[temp_w*6 +:temp_w] = v1428obus[temp_w*0 +:temp_w];
assign v1428ibus[data_w*0 +:data_w] = c180obus[data_w*6 +:data_w];
assign c181ibus[temp_w*0 +:temp_w] = v112obus[temp_w*1 +:temp_w];
assign v112ibus[data_w*1 +:data_w] = c181obus[data_w*0 +:data_w];
assign c181ibus[temp_w*1 +:temp_w] = v491obus[temp_w*0 +:temp_w];
assign v491ibus[data_w*0 +:data_w] = c181obus[data_w*1 +:data_w];
assign c181ibus[temp_w*2 +:temp_w] = v644obus[temp_w*0 +:temp_w];
assign v644ibus[data_w*0 +:data_w] = c181obus[data_w*2 +:data_w];
assign c181ibus[temp_w*3 +:temp_w] = v766obus[temp_w*0 +:temp_w];
assign v766ibus[data_w*0 +:data_w] = c181obus[data_w*3 +:data_w];
assign c181ibus[temp_w*4 +:temp_w] = v1057obus[temp_w*0 +:temp_w];
assign v1057ibus[data_w*0 +:data_w] = c181obus[data_w*4 +:data_w];
assign c181ibus[temp_w*5 +:temp_w] = v1333obus[temp_w*1 +:temp_w];
assign v1333ibus[data_w*1 +:data_w] = c181obus[data_w*5 +:data_w];
assign c181ibus[temp_w*6 +:temp_w] = v1429obus[temp_w*0 +:temp_w];
assign v1429ibus[data_w*0 +:data_w] = c181obus[data_w*6 +:data_w];
assign c182ibus[temp_w*0 +:temp_w] = v113obus[temp_w*1 +:temp_w];
assign v113ibus[data_w*1 +:data_w] = c182obus[data_w*0 +:data_w];
assign c182ibus[temp_w*1 +:temp_w] = v492obus[temp_w*0 +:temp_w];
assign v492ibus[data_w*0 +:data_w] = c182obus[data_w*1 +:data_w];
assign c182ibus[temp_w*2 +:temp_w] = v645obus[temp_w*0 +:temp_w];
assign v645ibus[data_w*0 +:data_w] = c182obus[data_w*2 +:data_w];
assign c182ibus[temp_w*3 +:temp_w] = v767obus[temp_w*0 +:temp_w];
assign v767ibus[data_w*0 +:data_w] = c182obus[data_w*3 +:data_w];
assign c182ibus[temp_w*4 +:temp_w] = v1058obus[temp_w*0 +:temp_w];
assign v1058ibus[data_w*0 +:data_w] = c182obus[data_w*4 +:data_w];
assign c182ibus[temp_w*5 +:temp_w] = v1334obus[temp_w*1 +:temp_w];
assign v1334ibus[data_w*1 +:data_w] = c182obus[data_w*5 +:data_w];
assign c182ibus[temp_w*6 +:temp_w] = v1430obus[temp_w*0 +:temp_w];
assign v1430ibus[data_w*0 +:data_w] = c182obus[data_w*6 +:data_w];
assign c183ibus[temp_w*0 +:temp_w] = v114obus[temp_w*1 +:temp_w];
assign v114ibus[data_w*1 +:data_w] = c183obus[data_w*0 +:data_w];
assign c183ibus[temp_w*1 +:temp_w] = v493obus[temp_w*0 +:temp_w];
assign v493ibus[data_w*0 +:data_w] = c183obus[data_w*1 +:data_w];
assign c183ibus[temp_w*2 +:temp_w] = v646obus[temp_w*0 +:temp_w];
assign v646ibus[data_w*0 +:data_w] = c183obus[data_w*2 +:data_w];
assign c183ibus[temp_w*3 +:temp_w] = v672obus[temp_w*0 +:temp_w];
assign v672ibus[data_w*0 +:data_w] = c183obus[data_w*3 +:data_w];
assign c183ibus[temp_w*4 +:temp_w] = v1059obus[temp_w*0 +:temp_w];
assign v1059ibus[data_w*0 +:data_w] = c183obus[data_w*4 +:data_w];
assign c183ibus[temp_w*5 +:temp_w] = v1335obus[temp_w*1 +:temp_w];
assign v1335ibus[data_w*1 +:data_w] = c183obus[data_w*5 +:data_w];
assign c183ibus[temp_w*6 +:temp_w] = v1431obus[temp_w*0 +:temp_w];
assign v1431ibus[data_w*0 +:data_w] = c183obus[data_w*6 +:data_w];
assign c184ibus[temp_w*0 +:temp_w] = v115obus[temp_w*1 +:temp_w];
assign v115ibus[data_w*1 +:data_w] = c184obus[data_w*0 +:data_w];
assign c184ibus[temp_w*1 +:temp_w] = v494obus[temp_w*0 +:temp_w];
assign v494ibus[data_w*0 +:data_w] = c184obus[data_w*1 +:data_w];
assign c184ibus[temp_w*2 +:temp_w] = v647obus[temp_w*0 +:temp_w];
assign v647ibus[data_w*0 +:data_w] = c184obus[data_w*2 +:data_w];
assign c184ibus[temp_w*3 +:temp_w] = v673obus[temp_w*0 +:temp_w];
assign v673ibus[data_w*0 +:data_w] = c184obus[data_w*3 +:data_w];
assign c184ibus[temp_w*4 +:temp_w] = v1060obus[temp_w*0 +:temp_w];
assign v1060ibus[data_w*0 +:data_w] = c184obus[data_w*4 +:data_w];
assign c184ibus[temp_w*5 +:temp_w] = v1336obus[temp_w*1 +:temp_w];
assign v1336ibus[data_w*1 +:data_w] = c184obus[data_w*5 +:data_w];
assign c184ibus[temp_w*6 +:temp_w] = v1432obus[temp_w*0 +:temp_w];
assign v1432ibus[data_w*0 +:data_w] = c184obus[data_w*6 +:data_w];
assign c185ibus[temp_w*0 +:temp_w] = v116obus[temp_w*1 +:temp_w];
assign v116ibus[data_w*1 +:data_w] = c185obus[data_w*0 +:data_w];
assign c185ibus[temp_w*1 +:temp_w] = v495obus[temp_w*0 +:temp_w];
assign v495ibus[data_w*0 +:data_w] = c185obus[data_w*1 +:data_w];
assign c185ibus[temp_w*2 +:temp_w] = v648obus[temp_w*0 +:temp_w];
assign v648ibus[data_w*0 +:data_w] = c185obus[data_w*2 +:data_w];
assign c185ibus[temp_w*3 +:temp_w] = v674obus[temp_w*0 +:temp_w];
assign v674ibus[data_w*0 +:data_w] = c185obus[data_w*3 +:data_w];
assign c185ibus[temp_w*4 +:temp_w] = v1061obus[temp_w*0 +:temp_w];
assign v1061ibus[data_w*0 +:data_w] = c185obus[data_w*4 +:data_w];
assign c185ibus[temp_w*5 +:temp_w] = v1337obus[temp_w*1 +:temp_w];
assign v1337ibus[data_w*1 +:data_w] = c185obus[data_w*5 +:data_w];
assign c185ibus[temp_w*6 +:temp_w] = v1433obus[temp_w*0 +:temp_w];
assign v1433ibus[data_w*0 +:data_w] = c185obus[data_w*6 +:data_w];
assign c186ibus[temp_w*0 +:temp_w] = v117obus[temp_w*1 +:temp_w];
assign v117ibus[data_w*1 +:data_w] = c186obus[data_w*0 +:data_w];
assign c186ibus[temp_w*1 +:temp_w] = v496obus[temp_w*0 +:temp_w];
assign v496ibus[data_w*0 +:data_w] = c186obus[data_w*1 +:data_w];
assign c186ibus[temp_w*2 +:temp_w] = v649obus[temp_w*0 +:temp_w];
assign v649ibus[data_w*0 +:data_w] = c186obus[data_w*2 +:data_w];
assign c186ibus[temp_w*3 +:temp_w] = v675obus[temp_w*0 +:temp_w];
assign v675ibus[data_w*0 +:data_w] = c186obus[data_w*3 +:data_w];
assign c186ibus[temp_w*4 +:temp_w] = v1062obus[temp_w*0 +:temp_w];
assign v1062ibus[data_w*0 +:data_w] = c186obus[data_w*4 +:data_w];
assign c186ibus[temp_w*5 +:temp_w] = v1338obus[temp_w*1 +:temp_w];
assign v1338ibus[data_w*1 +:data_w] = c186obus[data_w*5 +:data_w];
assign c186ibus[temp_w*6 +:temp_w] = v1434obus[temp_w*0 +:temp_w];
assign v1434ibus[data_w*0 +:data_w] = c186obus[data_w*6 +:data_w];
assign c187ibus[temp_w*0 +:temp_w] = v118obus[temp_w*1 +:temp_w];
assign v118ibus[data_w*1 +:data_w] = c187obus[data_w*0 +:data_w];
assign c187ibus[temp_w*1 +:temp_w] = v497obus[temp_w*0 +:temp_w];
assign v497ibus[data_w*0 +:data_w] = c187obus[data_w*1 +:data_w];
assign c187ibus[temp_w*2 +:temp_w] = v650obus[temp_w*0 +:temp_w];
assign v650ibus[data_w*0 +:data_w] = c187obus[data_w*2 +:data_w];
assign c187ibus[temp_w*3 +:temp_w] = v676obus[temp_w*0 +:temp_w];
assign v676ibus[data_w*0 +:data_w] = c187obus[data_w*3 +:data_w];
assign c187ibus[temp_w*4 +:temp_w] = v1063obus[temp_w*0 +:temp_w];
assign v1063ibus[data_w*0 +:data_w] = c187obus[data_w*4 +:data_w];
assign c187ibus[temp_w*5 +:temp_w] = v1339obus[temp_w*1 +:temp_w];
assign v1339ibus[data_w*1 +:data_w] = c187obus[data_w*5 +:data_w];
assign c187ibus[temp_w*6 +:temp_w] = v1435obus[temp_w*0 +:temp_w];
assign v1435ibus[data_w*0 +:data_w] = c187obus[data_w*6 +:data_w];
assign c188ibus[temp_w*0 +:temp_w] = v119obus[temp_w*1 +:temp_w];
assign v119ibus[data_w*1 +:data_w] = c188obus[data_w*0 +:data_w];
assign c188ibus[temp_w*1 +:temp_w] = v498obus[temp_w*0 +:temp_w];
assign v498ibus[data_w*0 +:data_w] = c188obus[data_w*1 +:data_w];
assign c188ibus[temp_w*2 +:temp_w] = v651obus[temp_w*0 +:temp_w];
assign v651ibus[data_w*0 +:data_w] = c188obus[data_w*2 +:data_w];
assign c188ibus[temp_w*3 +:temp_w] = v677obus[temp_w*0 +:temp_w];
assign v677ibus[data_w*0 +:data_w] = c188obus[data_w*3 +:data_w];
assign c188ibus[temp_w*4 +:temp_w] = v1064obus[temp_w*0 +:temp_w];
assign v1064ibus[data_w*0 +:data_w] = c188obus[data_w*4 +:data_w];
assign c188ibus[temp_w*5 +:temp_w] = v1340obus[temp_w*1 +:temp_w];
assign v1340ibus[data_w*1 +:data_w] = c188obus[data_w*5 +:data_w];
assign c188ibus[temp_w*6 +:temp_w] = v1436obus[temp_w*0 +:temp_w];
assign v1436ibus[data_w*0 +:data_w] = c188obus[data_w*6 +:data_w];
assign c189ibus[temp_w*0 +:temp_w] = v120obus[temp_w*1 +:temp_w];
assign v120ibus[data_w*1 +:data_w] = c189obus[data_w*0 +:data_w];
assign c189ibus[temp_w*1 +:temp_w] = v499obus[temp_w*0 +:temp_w];
assign v499ibus[data_w*0 +:data_w] = c189obus[data_w*1 +:data_w];
assign c189ibus[temp_w*2 +:temp_w] = v652obus[temp_w*0 +:temp_w];
assign v652ibus[data_w*0 +:data_w] = c189obus[data_w*2 +:data_w];
assign c189ibus[temp_w*3 +:temp_w] = v678obus[temp_w*0 +:temp_w];
assign v678ibus[data_w*0 +:data_w] = c189obus[data_w*3 +:data_w];
assign c189ibus[temp_w*4 +:temp_w] = v1065obus[temp_w*0 +:temp_w];
assign v1065ibus[data_w*0 +:data_w] = c189obus[data_w*4 +:data_w];
assign c189ibus[temp_w*5 +:temp_w] = v1341obus[temp_w*1 +:temp_w];
assign v1341ibus[data_w*1 +:data_w] = c189obus[data_w*5 +:data_w];
assign c189ibus[temp_w*6 +:temp_w] = v1437obus[temp_w*0 +:temp_w];
assign v1437ibus[data_w*0 +:data_w] = c189obus[data_w*6 +:data_w];
assign c190ibus[temp_w*0 +:temp_w] = v121obus[temp_w*1 +:temp_w];
assign v121ibus[data_w*1 +:data_w] = c190obus[data_w*0 +:data_w];
assign c190ibus[temp_w*1 +:temp_w] = v500obus[temp_w*0 +:temp_w];
assign v500ibus[data_w*0 +:data_w] = c190obus[data_w*1 +:data_w];
assign c190ibus[temp_w*2 +:temp_w] = v653obus[temp_w*0 +:temp_w];
assign v653ibus[data_w*0 +:data_w] = c190obus[data_w*2 +:data_w];
assign c190ibus[temp_w*3 +:temp_w] = v679obus[temp_w*0 +:temp_w];
assign v679ibus[data_w*0 +:data_w] = c190obus[data_w*3 +:data_w];
assign c190ibus[temp_w*4 +:temp_w] = v1066obus[temp_w*0 +:temp_w];
assign v1066ibus[data_w*0 +:data_w] = c190obus[data_w*4 +:data_w];
assign c190ibus[temp_w*5 +:temp_w] = v1342obus[temp_w*1 +:temp_w];
assign v1342ibus[data_w*1 +:data_w] = c190obus[data_w*5 +:data_w];
assign c190ibus[temp_w*6 +:temp_w] = v1438obus[temp_w*0 +:temp_w];
assign v1438ibus[data_w*0 +:data_w] = c190obus[data_w*6 +:data_w];
assign c191ibus[temp_w*0 +:temp_w] = v122obus[temp_w*1 +:temp_w];
assign v122ibus[data_w*1 +:data_w] = c191obus[data_w*0 +:data_w];
assign c191ibus[temp_w*1 +:temp_w] = v501obus[temp_w*0 +:temp_w];
assign v501ibus[data_w*0 +:data_w] = c191obus[data_w*1 +:data_w];
assign c191ibus[temp_w*2 +:temp_w] = v654obus[temp_w*0 +:temp_w];
assign v654ibus[data_w*0 +:data_w] = c191obus[data_w*2 +:data_w];
assign c191ibus[temp_w*3 +:temp_w] = v680obus[temp_w*0 +:temp_w];
assign v680ibus[data_w*0 +:data_w] = c191obus[data_w*3 +:data_w];
assign c191ibus[temp_w*4 +:temp_w] = v1067obus[temp_w*0 +:temp_w];
assign v1067ibus[data_w*0 +:data_w] = c191obus[data_w*4 +:data_w];
assign c191ibus[temp_w*5 +:temp_w] = v1343obus[temp_w*1 +:temp_w];
assign v1343ibus[data_w*1 +:data_w] = c191obus[data_w*5 +:data_w];
assign c191ibus[temp_w*6 +:temp_w] = v1439obus[temp_w*0 +:temp_w];
assign v1439ibus[data_w*0 +:data_w] = c191obus[data_w*6 +:data_w];
assign c192ibus[temp_w*0 +:temp_w] = v312obus[temp_w*0 +:temp_w];
assign v312ibus[data_w*0 +:data_w] = c192obus[data_w*0 +:data_w];
assign c192ibus[temp_w*1 +:temp_w] = v406obus[temp_w*0 +:temp_w];
assign v406ibus[data_w*0 +:data_w] = c192obus[data_w*1 +:data_w];
assign c192ibus[temp_w*2 +:temp_w] = v561obus[temp_w*1 +:temp_w];
assign v561ibus[data_w*1 +:data_w] = c192obus[data_w*2 +:data_w];
assign c192ibus[temp_w*3 +:temp_w] = v705obus[temp_w*1 +:temp_w];
assign v705ibus[data_w*1 +:data_w] = c192obus[data_w*3 +:data_w];
assign c192ibus[temp_w*4 +:temp_w] = v1056obus[temp_w*1 +:temp_w];
assign v1056ibus[data_w*1 +:data_w] = c192obus[data_w*4 +:data_w];
assign c192ibus[temp_w*5 +:temp_w] = v1344obus[temp_w*1 +:temp_w];
assign v1344ibus[data_w*1 +:data_w] = c192obus[data_w*5 +:data_w];
assign c192ibus[temp_w*6 +:temp_w] = v1440obus[temp_w*0 +:temp_w];
assign v1440ibus[data_w*0 +:data_w] = c192obus[data_w*6 +:data_w];
assign c193ibus[temp_w*0 +:temp_w] = v313obus[temp_w*0 +:temp_w];
assign v313ibus[data_w*0 +:data_w] = c193obus[data_w*0 +:data_w];
assign c193ibus[temp_w*1 +:temp_w] = v407obus[temp_w*0 +:temp_w];
assign v407ibus[data_w*0 +:data_w] = c193obus[data_w*1 +:data_w];
assign c193ibus[temp_w*2 +:temp_w] = v562obus[temp_w*1 +:temp_w];
assign v562ibus[data_w*1 +:data_w] = c193obus[data_w*2 +:data_w];
assign c193ibus[temp_w*3 +:temp_w] = v706obus[temp_w*1 +:temp_w];
assign v706ibus[data_w*1 +:data_w] = c193obus[data_w*3 +:data_w];
assign c193ibus[temp_w*4 +:temp_w] = v1057obus[temp_w*1 +:temp_w];
assign v1057ibus[data_w*1 +:data_w] = c193obus[data_w*4 +:data_w];
assign c193ibus[temp_w*5 +:temp_w] = v1345obus[temp_w*1 +:temp_w];
assign v1345ibus[data_w*1 +:data_w] = c193obus[data_w*5 +:data_w];
assign c193ibus[temp_w*6 +:temp_w] = v1441obus[temp_w*0 +:temp_w];
assign v1441ibus[data_w*0 +:data_w] = c193obus[data_w*6 +:data_w];
assign c194ibus[temp_w*0 +:temp_w] = v314obus[temp_w*0 +:temp_w];
assign v314ibus[data_w*0 +:data_w] = c194obus[data_w*0 +:data_w];
assign c194ibus[temp_w*1 +:temp_w] = v408obus[temp_w*0 +:temp_w];
assign v408ibus[data_w*0 +:data_w] = c194obus[data_w*1 +:data_w];
assign c194ibus[temp_w*2 +:temp_w] = v563obus[temp_w*1 +:temp_w];
assign v563ibus[data_w*1 +:data_w] = c194obus[data_w*2 +:data_w];
assign c194ibus[temp_w*3 +:temp_w] = v707obus[temp_w*1 +:temp_w];
assign v707ibus[data_w*1 +:data_w] = c194obus[data_w*3 +:data_w];
assign c194ibus[temp_w*4 +:temp_w] = v1058obus[temp_w*1 +:temp_w];
assign v1058ibus[data_w*1 +:data_w] = c194obus[data_w*4 +:data_w];
assign c194ibus[temp_w*5 +:temp_w] = v1346obus[temp_w*1 +:temp_w];
assign v1346ibus[data_w*1 +:data_w] = c194obus[data_w*5 +:data_w];
assign c194ibus[temp_w*6 +:temp_w] = v1442obus[temp_w*0 +:temp_w];
assign v1442ibus[data_w*0 +:data_w] = c194obus[data_w*6 +:data_w];
assign c195ibus[temp_w*0 +:temp_w] = v315obus[temp_w*0 +:temp_w];
assign v315ibus[data_w*0 +:data_w] = c195obus[data_w*0 +:data_w];
assign c195ibus[temp_w*1 +:temp_w] = v409obus[temp_w*0 +:temp_w];
assign v409ibus[data_w*0 +:data_w] = c195obus[data_w*1 +:data_w];
assign c195ibus[temp_w*2 +:temp_w] = v564obus[temp_w*1 +:temp_w];
assign v564ibus[data_w*1 +:data_w] = c195obus[data_w*2 +:data_w];
assign c195ibus[temp_w*3 +:temp_w] = v708obus[temp_w*1 +:temp_w];
assign v708ibus[data_w*1 +:data_w] = c195obus[data_w*3 +:data_w];
assign c195ibus[temp_w*4 +:temp_w] = v1059obus[temp_w*1 +:temp_w];
assign v1059ibus[data_w*1 +:data_w] = c195obus[data_w*4 +:data_w];
assign c195ibus[temp_w*5 +:temp_w] = v1347obus[temp_w*1 +:temp_w];
assign v1347ibus[data_w*1 +:data_w] = c195obus[data_w*5 +:data_w];
assign c195ibus[temp_w*6 +:temp_w] = v1443obus[temp_w*0 +:temp_w];
assign v1443ibus[data_w*0 +:data_w] = c195obus[data_w*6 +:data_w];
assign c196ibus[temp_w*0 +:temp_w] = v316obus[temp_w*0 +:temp_w];
assign v316ibus[data_w*0 +:data_w] = c196obus[data_w*0 +:data_w];
assign c196ibus[temp_w*1 +:temp_w] = v410obus[temp_w*0 +:temp_w];
assign v410ibus[data_w*0 +:data_w] = c196obus[data_w*1 +:data_w];
assign c196ibus[temp_w*2 +:temp_w] = v565obus[temp_w*1 +:temp_w];
assign v565ibus[data_w*1 +:data_w] = c196obus[data_w*2 +:data_w];
assign c196ibus[temp_w*3 +:temp_w] = v709obus[temp_w*1 +:temp_w];
assign v709ibus[data_w*1 +:data_w] = c196obus[data_w*3 +:data_w];
assign c196ibus[temp_w*4 +:temp_w] = v1060obus[temp_w*1 +:temp_w];
assign v1060ibus[data_w*1 +:data_w] = c196obus[data_w*4 +:data_w];
assign c196ibus[temp_w*5 +:temp_w] = v1348obus[temp_w*1 +:temp_w];
assign v1348ibus[data_w*1 +:data_w] = c196obus[data_w*5 +:data_w];
assign c196ibus[temp_w*6 +:temp_w] = v1444obus[temp_w*0 +:temp_w];
assign v1444ibus[data_w*0 +:data_w] = c196obus[data_w*6 +:data_w];
assign c197ibus[temp_w*0 +:temp_w] = v317obus[temp_w*0 +:temp_w];
assign v317ibus[data_w*0 +:data_w] = c197obus[data_w*0 +:data_w];
assign c197ibus[temp_w*1 +:temp_w] = v411obus[temp_w*0 +:temp_w];
assign v411ibus[data_w*0 +:data_w] = c197obus[data_w*1 +:data_w];
assign c197ibus[temp_w*2 +:temp_w] = v566obus[temp_w*1 +:temp_w];
assign v566ibus[data_w*1 +:data_w] = c197obus[data_w*2 +:data_w];
assign c197ibus[temp_w*3 +:temp_w] = v710obus[temp_w*1 +:temp_w];
assign v710ibus[data_w*1 +:data_w] = c197obus[data_w*3 +:data_w];
assign c197ibus[temp_w*4 +:temp_w] = v1061obus[temp_w*1 +:temp_w];
assign v1061ibus[data_w*1 +:data_w] = c197obus[data_w*4 +:data_w];
assign c197ibus[temp_w*5 +:temp_w] = v1349obus[temp_w*1 +:temp_w];
assign v1349ibus[data_w*1 +:data_w] = c197obus[data_w*5 +:data_w];
assign c197ibus[temp_w*6 +:temp_w] = v1445obus[temp_w*0 +:temp_w];
assign v1445ibus[data_w*0 +:data_w] = c197obus[data_w*6 +:data_w];
assign c198ibus[temp_w*0 +:temp_w] = v318obus[temp_w*0 +:temp_w];
assign v318ibus[data_w*0 +:data_w] = c198obus[data_w*0 +:data_w];
assign c198ibus[temp_w*1 +:temp_w] = v412obus[temp_w*0 +:temp_w];
assign v412ibus[data_w*0 +:data_w] = c198obus[data_w*1 +:data_w];
assign c198ibus[temp_w*2 +:temp_w] = v567obus[temp_w*1 +:temp_w];
assign v567ibus[data_w*1 +:data_w] = c198obus[data_w*2 +:data_w];
assign c198ibus[temp_w*3 +:temp_w] = v711obus[temp_w*1 +:temp_w];
assign v711ibus[data_w*1 +:data_w] = c198obus[data_w*3 +:data_w];
assign c198ibus[temp_w*4 +:temp_w] = v1062obus[temp_w*1 +:temp_w];
assign v1062ibus[data_w*1 +:data_w] = c198obus[data_w*4 +:data_w];
assign c198ibus[temp_w*5 +:temp_w] = v1350obus[temp_w*1 +:temp_w];
assign v1350ibus[data_w*1 +:data_w] = c198obus[data_w*5 +:data_w];
assign c198ibus[temp_w*6 +:temp_w] = v1446obus[temp_w*0 +:temp_w];
assign v1446ibus[data_w*0 +:data_w] = c198obus[data_w*6 +:data_w];
assign c199ibus[temp_w*0 +:temp_w] = v319obus[temp_w*0 +:temp_w];
assign v319ibus[data_w*0 +:data_w] = c199obus[data_w*0 +:data_w];
assign c199ibus[temp_w*1 +:temp_w] = v413obus[temp_w*0 +:temp_w];
assign v413ibus[data_w*0 +:data_w] = c199obus[data_w*1 +:data_w];
assign c199ibus[temp_w*2 +:temp_w] = v568obus[temp_w*1 +:temp_w];
assign v568ibus[data_w*1 +:data_w] = c199obus[data_w*2 +:data_w];
assign c199ibus[temp_w*3 +:temp_w] = v712obus[temp_w*1 +:temp_w];
assign v712ibus[data_w*1 +:data_w] = c199obus[data_w*3 +:data_w];
assign c199ibus[temp_w*4 +:temp_w] = v1063obus[temp_w*1 +:temp_w];
assign v1063ibus[data_w*1 +:data_w] = c199obus[data_w*4 +:data_w];
assign c199ibus[temp_w*5 +:temp_w] = v1351obus[temp_w*1 +:temp_w];
assign v1351ibus[data_w*1 +:data_w] = c199obus[data_w*5 +:data_w];
assign c199ibus[temp_w*6 +:temp_w] = v1447obus[temp_w*0 +:temp_w];
assign v1447ibus[data_w*0 +:data_w] = c199obus[data_w*6 +:data_w];
assign c200ibus[temp_w*0 +:temp_w] = v320obus[temp_w*0 +:temp_w];
assign v320ibus[data_w*0 +:data_w] = c200obus[data_w*0 +:data_w];
assign c200ibus[temp_w*1 +:temp_w] = v414obus[temp_w*0 +:temp_w];
assign v414ibus[data_w*0 +:data_w] = c200obus[data_w*1 +:data_w];
assign c200ibus[temp_w*2 +:temp_w] = v569obus[temp_w*1 +:temp_w];
assign v569ibus[data_w*1 +:data_w] = c200obus[data_w*2 +:data_w];
assign c200ibus[temp_w*3 +:temp_w] = v713obus[temp_w*1 +:temp_w];
assign v713ibus[data_w*1 +:data_w] = c200obus[data_w*3 +:data_w];
assign c200ibus[temp_w*4 +:temp_w] = v1064obus[temp_w*1 +:temp_w];
assign v1064ibus[data_w*1 +:data_w] = c200obus[data_w*4 +:data_w];
assign c200ibus[temp_w*5 +:temp_w] = v1352obus[temp_w*1 +:temp_w];
assign v1352ibus[data_w*1 +:data_w] = c200obus[data_w*5 +:data_w];
assign c200ibus[temp_w*6 +:temp_w] = v1448obus[temp_w*0 +:temp_w];
assign v1448ibus[data_w*0 +:data_w] = c200obus[data_w*6 +:data_w];
assign c201ibus[temp_w*0 +:temp_w] = v321obus[temp_w*0 +:temp_w];
assign v321ibus[data_w*0 +:data_w] = c201obus[data_w*0 +:data_w];
assign c201ibus[temp_w*1 +:temp_w] = v415obus[temp_w*0 +:temp_w];
assign v415ibus[data_w*0 +:data_w] = c201obus[data_w*1 +:data_w];
assign c201ibus[temp_w*2 +:temp_w] = v570obus[temp_w*1 +:temp_w];
assign v570ibus[data_w*1 +:data_w] = c201obus[data_w*2 +:data_w];
assign c201ibus[temp_w*3 +:temp_w] = v714obus[temp_w*1 +:temp_w];
assign v714ibus[data_w*1 +:data_w] = c201obus[data_w*3 +:data_w];
assign c201ibus[temp_w*4 +:temp_w] = v1065obus[temp_w*1 +:temp_w];
assign v1065ibus[data_w*1 +:data_w] = c201obus[data_w*4 +:data_w];
assign c201ibus[temp_w*5 +:temp_w] = v1353obus[temp_w*1 +:temp_w];
assign v1353ibus[data_w*1 +:data_w] = c201obus[data_w*5 +:data_w];
assign c201ibus[temp_w*6 +:temp_w] = v1449obus[temp_w*0 +:temp_w];
assign v1449ibus[data_w*0 +:data_w] = c201obus[data_w*6 +:data_w];
assign c202ibus[temp_w*0 +:temp_w] = v322obus[temp_w*0 +:temp_w];
assign v322ibus[data_w*0 +:data_w] = c202obus[data_w*0 +:data_w];
assign c202ibus[temp_w*1 +:temp_w] = v416obus[temp_w*0 +:temp_w];
assign v416ibus[data_w*0 +:data_w] = c202obus[data_w*1 +:data_w];
assign c202ibus[temp_w*2 +:temp_w] = v571obus[temp_w*1 +:temp_w];
assign v571ibus[data_w*1 +:data_w] = c202obus[data_w*2 +:data_w];
assign c202ibus[temp_w*3 +:temp_w] = v715obus[temp_w*1 +:temp_w];
assign v715ibus[data_w*1 +:data_w] = c202obus[data_w*3 +:data_w];
assign c202ibus[temp_w*4 +:temp_w] = v1066obus[temp_w*1 +:temp_w];
assign v1066ibus[data_w*1 +:data_w] = c202obus[data_w*4 +:data_w];
assign c202ibus[temp_w*5 +:temp_w] = v1354obus[temp_w*1 +:temp_w];
assign v1354ibus[data_w*1 +:data_w] = c202obus[data_w*5 +:data_w];
assign c202ibus[temp_w*6 +:temp_w] = v1450obus[temp_w*0 +:temp_w];
assign v1450ibus[data_w*0 +:data_w] = c202obus[data_w*6 +:data_w];
assign c203ibus[temp_w*0 +:temp_w] = v323obus[temp_w*0 +:temp_w];
assign v323ibus[data_w*0 +:data_w] = c203obus[data_w*0 +:data_w];
assign c203ibus[temp_w*1 +:temp_w] = v417obus[temp_w*0 +:temp_w];
assign v417ibus[data_w*0 +:data_w] = c203obus[data_w*1 +:data_w];
assign c203ibus[temp_w*2 +:temp_w] = v572obus[temp_w*1 +:temp_w];
assign v572ibus[data_w*1 +:data_w] = c203obus[data_w*2 +:data_w];
assign c203ibus[temp_w*3 +:temp_w] = v716obus[temp_w*1 +:temp_w];
assign v716ibus[data_w*1 +:data_w] = c203obus[data_w*3 +:data_w];
assign c203ibus[temp_w*4 +:temp_w] = v1067obus[temp_w*1 +:temp_w];
assign v1067ibus[data_w*1 +:data_w] = c203obus[data_w*4 +:data_w];
assign c203ibus[temp_w*5 +:temp_w] = v1355obus[temp_w*1 +:temp_w];
assign v1355ibus[data_w*1 +:data_w] = c203obus[data_w*5 +:data_w];
assign c203ibus[temp_w*6 +:temp_w] = v1451obus[temp_w*0 +:temp_w];
assign v1451ibus[data_w*0 +:data_w] = c203obus[data_w*6 +:data_w];
assign c204ibus[temp_w*0 +:temp_w] = v324obus[temp_w*0 +:temp_w];
assign v324ibus[data_w*0 +:data_w] = c204obus[data_w*0 +:data_w];
assign c204ibus[temp_w*1 +:temp_w] = v418obus[temp_w*0 +:temp_w];
assign v418ibus[data_w*0 +:data_w] = c204obus[data_w*1 +:data_w];
assign c204ibus[temp_w*2 +:temp_w] = v573obus[temp_w*1 +:temp_w];
assign v573ibus[data_w*1 +:data_w] = c204obus[data_w*2 +:data_w];
assign c204ibus[temp_w*3 +:temp_w] = v717obus[temp_w*1 +:temp_w];
assign v717ibus[data_w*1 +:data_w] = c204obus[data_w*3 +:data_w];
assign c204ibus[temp_w*4 +:temp_w] = v1068obus[temp_w*1 +:temp_w];
assign v1068ibus[data_w*1 +:data_w] = c204obus[data_w*4 +:data_w];
assign c204ibus[temp_w*5 +:temp_w] = v1356obus[temp_w*1 +:temp_w];
assign v1356ibus[data_w*1 +:data_w] = c204obus[data_w*5 +:data_w];
assign c204ibus[temp_w*6 +:temp_w] = v1452obus[temp_w*0 +:temp_w];
assign v1452ibus[data_w*0 +:data_w] = c204obus[data_w*6 +:data_w];
assign c205ibus[temp_w*0 +:temp_w] = v325obus[temp_w*0 +:temp_w];
assign v325ibus[data_w*0 +:data_w] = c205obus[data_w*0 +:data_w];
assign c205ibus[temp_w*1 +:temp_w] = v419obus[temp_w*0 +:temp_w];
assign v419ibus[data_w*0 +:data_w] = c205obus[data_w*1 +:data_w];
assign c205ibus[temp_w*2 +:temp_w] = v574obus[temp_w*1 +:temp_w];
assign v574ibus[data_w*1 +:data_w] = c205obus[data_w*2 +:data_w];
assign c205ibus[temp_w*3 +:temp_w] = v718obus[temp_w*1 +:temp_w];
assign v718ibus[data_w*1 +:data_w] = c205obus[data_w*3 +:data_w];
assign c205ibus[temp_w*4 +:temp_w] = v1069obus[temp_w*1 +:temp_w];
assign v1069ibus[data_w*1 +:data_w] = c205obus[data_w*4 +:data_w];
assign c205ibus[temp_w*5 +:temp_w] = v1357obus[temp_w*1 +:temp_w];
assign v1357ibus[data_w*1 +:data_w] = c205obus[data_w*5 +:data_w];
assign c205ibus[temp_w*6 +:temp_w] = v1453obus[temp_w*0 +:temp_w];
assign v1453ibus[data_w*0 +:data_w] = c205obus[data_w*6 +:data_w];
assign c206ibus[temp_w*0 +:temp_w] = v326obus[temp_w*0 +:temp_w];
assign v326ibus[data_w*0 +:data_w] = c206obus[data_w*0 +:data_w];
assign c206ibus[temp_w*1 +:temp_w] = v420obus[temp_w*0 +:temp_w];
assign v420ibus[data_w*0 +:data_w] = c206obus[data_w*1 +:data_w];
assign c206ibus[temp_w*2 +:temp_w] = v575obus[temp_w*1 +:temp_w];
assign v575ibus[data_w*1 +:data_w] = c206obus[data_w*2 +:data_w];
assign c206ibus[temp_w*3 +:temp_w] = v719obus[temp_w*1 +:temp_w];
assign v719ibus[data_w*1 +:data_w] = c206obus[data_w*3 +:data_w];
assign c206ibus[temp_w*4 +:temp_w] = v1070obus[temp_w*1 +:temp_w];
assign v1070ibus[data_w*1 +:data_w] = c206obus[data_w*4 +:data_w];
assign c206ibus[temp_w*5 +:temp_w] = v1358obus[temp_w*1 +:temp_w];
assign v1358ibus[data_w*1 +:data_w] = c206obus[data_w*5 +:data_w];
assign c206ibus[temp_w*6 +:temp_w] = v1454obus[temp_w*0 +:temp_w];
assign v1454ibus[data_w*0 +:data_w] = c206obus[data_w*6 +:data_w];
assign c207ibus[temp_w*0 +:temp_w] = v327obus[temp_w*0 +:temp_w];
assign v327ibus[data_w*0 +:data_w] = c207obus[data_w*0 +:data_w];
assign c207ibus[temp_w*1 +:temp_w] = v421obus[temp_w*0 +:temp_w];
assign v421ibus[data_w*0 +:data_w] = c207obus[data_w*1 +:data_w];
assign c207ibus[temp_w*2 +:temp_w] = v480obus[temp_w*1 +:temp_w];
assign v480ibus[data_w*1 +:data_w] = c207obus[data_w*2 +:data_w];
assign c207ibus[temp_w*3 +:temp_w] = v720obus[temp_w*1 +:temp_w];
assign v720ibus[data_w*1 +:data_w] = c207obus[data_w*3 +:data_w];
assign c207ibus[temp_w*4 +:temp_w] = v1071obus[temp_w*1 +:temp_w];
assign v1071ibus[data_w*1 +:data_w] = c207obus[data_w*4 +:data_w];
assign c207ibus[temp_w*5 +:temp_w] = v1359obus[temp_w*1 +:temp_w];
assign v1359ibus[data_w*1 +:data_w] = c207obus[data_w*5 +:data_w];
assign c207ibus[temp_w*6 +:temp_w] = v1455obus[temp_w*0 +:temp_w];
assign v1455ibus[data_w*0 +:data_w] = c207obus[data_w*6 +:data_w];
assign c208ibus[temp_w*0 +:temp_w] = v328obus[temp_w*0 +:temp_w];
assign v328ibus[data_w*0 +:data_w] = c208obus[data_w*0 +:data_w];
assign c208ibus[temp_w*1 +:temp_w] = v422obus[temp_w*0 +:temp_w];
assign v422ibus[data_w*0 +:data_w] = c208obus[data_w*1 +:data_w];
assign c208ibus[temp_w*2 +:temp_w] = v481obus[temp_w*1 +:temp_w];
assign v481ibus[data_w*1 +:data_w] = c208obus[data_w*2 +:data_w];
assign c208ibus[temp_w*3 +:temp_w] = v721obus[temp_w*1 +:temp_w];
assign v721ibus[data_w*1 +:data_w] = c208obus[data_w*3 +:data_w];
assign c208ibus[temp_w*4 +:temp_w] = v1072obus[temp_w*1 +:temp_w];
assign v1072ibus[data_w*1 +:data_w] = c208obus[data_w*4 +:data_w];
assign c208ibus[temp_w*5 +:temp_w] = v1360obus[temp_w*1 +:temp_w];
assign v1360ibus[data_w*1 +:data_w] = c208obus[data_w*5 +:data_w];
assign c208ibus[temp_w*6 +:temp_w] = v1456obus[temp_w*0 +:temp_w];
assign v1456ibus[data_w*0 +:data_w] = c208obus[data_w*6 +:data_w];
assign c209ibus[temp_w*0 +:temp_w] = v329obus[temp_w*0 +:temp_w];
assign v329ibus[data_w*0 +:data_w] = c209obus[data_w*0 +:data_w];
assign c209ibus[temp_w*1 +:temp_w] = v423obus[temp_w*0 +:temp_w];
assign v423ibus[data_w*0 +:data_w] = c209obus[data_w*1 +:data_w];
assign c209ibus[temp_w*2 +:temp_w] = v482obus[temp_w*1 +:temp_w];
assign v482ibus[data_w*1 +:data_w] = c209obus[data_w*2 +:data_w];
assign c209ibus[temp_w*3 +:temp_w] = v722obus[temp_w*1 +:temp_w];
assign v722ibus[data_w*1 +:data_w] = c209obus[data_w*3 +:data_w];
assign c209ibus[temp_w*4 +:temp_w] = v1073obus[temp_w*1 +:temp_w];
assign v1073ibus[data_w*1 +:data_w] = c209obus[data_w*4 +:data_w];
assign c209ibus[temp_w*5 +:temp_w] = v1361obus[temp_w*1 +:temp_w];
assign v1361ibus[data_w*1 +:data_w] = c209obus[data_w*5 +:data_w];
assign c209ibus[temp_w*6 +:temp_w] = v1457obus[temp_w*0 +:temp_w];
assign v1457ibus[data_w*0 +:data_w] = c209obus[data_w*6 +:data_w];
assign c210ibus[temp_w*0 +:temp_w] = v330obus[temp_w*0 +:temp_w];
assign v330ibus[data_w*0 +:data_w] = c210obus[data_w*0 +:data_w];
assign c210ibus[temp_w*1 +:temp_w] = v424obus[temp_w*0 +:temp_w];
assign v424ibus[data_w*0 +:data_w] = c210obus[data_w*1 +:data_w];
assign c210ibus[temp_w*2 +:temp_w] = v483obus[temp_w*1 +:temp_w];
assign v483ibus[data_w*1 +:data_w] = c210obus[data_w*2 +:data_w];
assign c210ibus[temp_w*3 +:temp_w] = v723obus[temp_w*1 +:temp_w];
assign v723ibus[data_w*1 +:data_w] = c210obus[data_w*3 +:data_w];
assign c210ibus[temp_w*4 +:temp_w] = v1074obus[temp_w*1 +:temp_w];
assign v1074ibus[data_w*1 +:data_w] = c210obus[data_w*4 +:data_w];
assign c210ibus[temp_w*5 +:temp_w] = v1362obus[temp_w*1 +:temp_w];
assign v1362ibus[data_w*1 +:data_w] = c210obus[data_w*5 +:data_w];
assign c210ibus[temp_w*6 +:temp_w] = v1458obus[temp_w*0 +:temp_w];
assign v1458ibus[data_w*0 +:data_w] = c210obus[data_w*6 +:data_w];
assign c211ibus[temp_w*0 +:temp_w] = v331obus[temp_w*0 +:temp_w];
assign v331ibus[data_w*0 +:data_w] = c211obus[data_w*0 +:data_w];
assign c211ibus[temp_w*1 +:temp_w] = v425obus[temp_w*0 +:temp_w];
assign v425ibus[data_w*0 +:data_w] = c211obus[data_w*1 +:data_w];
assign c211ibus[temp_w*2 +:temp_w] = v484obus[temp_w*1 +:temp_w];
assign v484ibus[data_w*1 +:data_w] = c211obus[data_w*2 +:data_w];
assign c211ibus[temp_w*3 +:temp_w] = v724obus[temp_w*1 +:temp_w];
assign v724ibus[data_w*1 +:data_w] = c211obus[data_w*3 +:data_w];
assign c211ibus[temp_w*4 +:temp_w] = v1075obus[temp_w*1 +:temp_w];
assign v1075ibus[data_w*1 +:data_w] = c211obus[data_w*4 +:data_w];
assign c211ibus[temp_w*5 +:temp_w] = v1363obus[temp_w*1 +:temp_w];
assign v1363ibus[data_w*1 +:data_w] = c211obus[data_w*5 +:data_w];
assign c211ibus[temp_w*6 +:temp_w] = v1459obus[temp_w*0 +:temp_w];
assign v1459ibus[data_w*0 +:data_w] = c211obus[data_w*6 +:data_w];
assign c212ibus[temp_w*0 +:temp_w] = v332obus[temp_w*0 +:temp_w];
assign v332ibus[data_w*0 +:data_w] = c212obus[data_w*0 +:data_w];
assign c212ibus[temp_w*1 +:temp_w] = v426obus[temp_w*0 +:temp_w];
assign v426ibus[data_w*0 +:data_w] = c212obus[data_w*1 +:data_w];
assign c212ibus[temp_w*2 +:temp_w] = v485obus[temp_w*1 +:temp_w];
assign v485ibus[data_w*1 +:data_w] = c212obus[data_w*2 +:data_w];
assign c212ibus[temp_w*3 +:temp_w] = v725obus[temp_w*1 +:temp_w];
assign v725ibus[data_w*1 +:data_w] = c212obus[data_w*3 +:data_w];
assign c212ibus[temp_w*4 +:temp_w] = v1076obus[temp_w*1 +:temp_w];
assign v1076ibus[data_w*1 +:data_w] = c212obus[data_w*4 +:data_w];
assign c212ibus[temp_w*5 +:temp_w] = v1364obus[temp_w*1 +:temp_w];
assign v1364ibus[data_w*1 +:data_w] = c212obus[data_w*5 +:data_w];
assign c212ibus[temp_w*6 +:temp_w] = v1460obus[temp_w*0 +:temp_w];
assign v1460ibus[data_w*0 +:data_w] = c212obus[data_w*6 +:data_w];
assign c213ibus[temp_w*0 +:temp_w] = v333obus[temp_w*0 +:temp_w];
assign v333ibus[data_w*0 +:data_w] = c213obus[data_w*0 +:data_w];
assign c213ibus[temp_w*1 +:temp_w] = v427obus[temp_w*0 +:temp_w];
assign v427ibus[data_w*0 +:data_w] = c213obus[data_w*1 +:data_w];
assign c213ibus[temp_w*2 +:temp_w] = v486obus[temp_w*1 +:temp_w];
assign v486ibus[data_w*1 +:data_w] = c213obus[data_w*2 +:data_w];
assign c213ibus[temp_w*3 +:temp_w] = v726obus[temp_w*1 +:temp_w];
assign v726ibus[data_w*1 +:data_w] = c213obus[data_w*3 +:data_w];
assign c213ibus[temp_w*4 +:temp_w] = v1077obus[temp_w*1 +:temp_w];
assign v1077ibus[data_w*1 +:data_w] = c213obus[data_w*4 +:data_w];
assign c213ibus[temp_w*5 +:temp_w] = v1365obus[temp_w*1 +:temp_w];
assign v1365ibus[data_w*1 +:data_w] = c213obus[data_w*5 +:data_w];
assign c213ibus[temp_w*6 +:temp_w] = v1461obus[temp_w*0 +:temp_w];
assign v1461ibus[data_w*0 +:data_w] = c213obus[data_w*6 +:data_w];
assign c214ibus[temp_w*0 +:temp_w] = v334obus[temp_w*0 +:temp_w];
assign v334ibus[data_w*0 +:data_w] = c214obus[data_w*0 +:data_w];
assign c214ibus[temp_w*1 +:temp_w] = v428obus[temp_w*0 +:temp_w];
assign v428ibus[data_w*0 +:data_w] = c214obus[data_w*1 +:data_w];
assign c214ibus[temp_w*2 +:temp_w] = v487obus[temp_w*1 +:temp_w];
assign v487ibus[data_w*1 +:data_w] = c214obus[data_w*2 +:data_w];
assign c214ibus[temp_w*3 +:temp_w] = v727obus[temp_w*1 +:temp_w];
assign v727ibus[data_w*1 +:data_w] = c214obus[data_w*3 +:data_w];
assign c214ibus[temp_w*4 +:temp_w] = v1078obus[temp_w*1 +:temp_w];
assign v1078ibus[data_w*1 +:data_w] = c214obus[data_w*4 +:data_w];
assign c214ibus[temp_w*5 +:temp_w] = v1366obus[temp_w*1 +:temp_w];
assign v1366ibus[data_w*1 +:data_w] = c214obus[data_w*5 +:data_w];
assign c214ibus[temp_w*6 +:temp_w] = v1462obus[temp_w*0 +:temp_w];
assign v1462ibus[data_w*0 +:data_w] = c214obus[data_w*6 +:data_w];
assign c215ibus[temp_w*0 +:temp_w] = v335obus[temp_w*0 +:temp_w];
assign v335ibus[data_w*0 +:data_w] = c215obus[data_w*0 +:data_w];
assign c215ibus[temp_w*1 +:temp_w] = v429obus[temp_w*0 +:temp_w];
assign v429ibus[data_w*0 +:data_w] = c215obus[data_w*1 +:data_w];
assign c215ibus[temp_w*2 +:temp_w] = v488obus[temp_w*1 +:temp_w];
assign v488ibus[data_w*1 +:data_w] = c215obus[data_w*2 +:data_w];
assign c215ibus[temp_w*3 +:temp_w] = v728obus[temp_w*1 +:temp_w];
assign v728ibus[data_w*1 +:data_w] = c215obus[data_w*3 +:data_w];
assign c215ibus[temp_w*4 +:temp_w] = v1079obus[temp_w*1 +:temp_w];
assign v1079ibus[data_w*1 +:data_w] = c215obus[data_w*4 +:data_w];
assign c215ibus[temp_w*5 +:temp_w] = v1367obus[temp_w*1 +:temp_w];
assign v1367ibus[data_w*1 +:data_w] = c215obus[data_w*5 +:data_w];
assign c215ibus[temp_w*6 +:temp_w] = v1463obus[temp_w*0 +:temp_w];
assign v1463ibus[data_w*0 +:data_w] = c215obus[data_w*6 +:data_w];
assign c216ibus[temp_w*0 +:temp_w] = v336obus[temp_w*0 +:temp_w];
assign v336ibus[data_w*0 +:data_w] = c216obus[data_w*0 +:data_w];
assign c216ibus[temp_w*1 +:temp_w] = v430obus[temp_w*0 +:temp_w];
assign v430ibus[data_w*0 +:data_w] = c216obus[data_w*1 +:data_w];
assign c216ibus[temp_w*2 +:temp_w] = v489obus[temp_w*1 +:temp_w];
assign v489ibus[data_w*1 +:data_w] = c216obus[data_w*2 +:data_w];
assign c216ibus[temp_w*3 +:temp_w] = v729obus[temp_w*1 +:temp_w];
assign v729ibus[data_w*1 +:data_w] = c216obus[data_w*3 +:data_w];
assign c216ibus[temp_w*4 +:temp_w] = v1080obus[temp_w*1 +:temp_w];
assign v1080ibus[data_w*1 +:data_w] = c216obus[data_w*4 +:data_w];
assign c216ibus[temp_w*5 +:temp_w] = v1368obus[temp_w*1 +:temp_w];
assign v1368ibus[data_w*1 +:data_w] = c216obus[data_w*5 +:data_w];
assign c216ibus[temp_w*6 +:temp_w] = v1464obus[temp_w*0 +:temp_w];
assign v1464ibus[data_w*0 +:data_w] = c216obus[data_w*6 +:data_w];
assign c217ibus[temp_w*0 +:temp_w] = v337obus[temp_w*0 +:temp_w];
assign v337ibus[data_w*0 +:data_w] = c217obus[data_w*0 +:data_w];
assign c217ibus[temp_w*1 +:temp_w] = v431obus[temp_w*0 +:temp_w];
assign v431ibus[data_w*0 +:data_w] = c217obus[data_w*1 +:data_w];
assign c217ibus[temp_w*2 +:temp_w] = v490obus[temp_w*1 +:temp_w];
assign v490ibus[data_w*1 +:data_w] = c217obus[data_w*2 +:data_w];
assign c217ibus[temp_w*3 +:temp_w] = v730obus[temp_w*1 +:temp_w];
assign v730ibus[data_w*1 +:data_w] = c217obus[data_w*3 +:data_w];
assign c217ibus[temp_w*4 +:temp_w] = v1081obus[temp_w*1 +:temp_w];
assign v1081ibus[data_w*1 +:data_w] = c217obus[data_w*4 +:data_w];
assign c217ibus[temp_w*5 +:temp_w] = v1369obus[temp_w*1 +:temp_w];
assign v1369ibus[data_w*1 +:data_w] = c217obus[data_w*5 +:data_w];
assign c217ibus[temp_w*6 +:temp_w] = v1465obus[temp_w*0 +:temp_w];
assign v1465ibus[data_w*0 +:data_w] = c217obus[data_w*6 +:data_w];
assign c218ibus[temp_w*0 +:temp_w] = v338obus[temp_w*0 +:temp_w];
assign v338ibus[data_w*0 +:data_w] = c218obus[data_w*0 +:data_w];
assign c218ibus[temp_w*1 +:temp_w] = v432obus[temp_w*0 +:temp_w];
assign v432ibus[data_w*0 +:data_w] = c218obus[data_w*1 +:data_w];
assign c218ibus[temp_w*2 +:temp_w] = v491obus[temp_w*1 +:temp_w];
assign v491ibus[data_w*1 +:data_w] = c218obus[data_w*2 +:data_w];
assign c218ibus[temp_w*3 +:temp_w] = v731obus[temp_w*1 +:temp_w];
assign v731ibus[data_w*1 +:data_w] = c218obus[data_w*3 +:data_w];
assign c218ibus[temp_w*4 +:temp_w] = v1082obus[temp_w*1 +:temp_w];
assign v1082ibus[data_w*1 +:data_w] = c218obus[data_w*4 +:data_w];
assign c218ibus[temp_w*5 +:temp_w] = v1370obus[temp_w*1 +:temp_w];
assign v1370ibus[data_w*1 +:data_w] = c218obus[data_w*5 +:data_w];
assign c218ibus[temp_w*6 +:temp_w] = v1466obus[temp_w*0 +:temp_w];
assign v1466ibus[data_w*0 +:data_w] = c218obus[data_w*6 +:data_w];
assign c219ibus[temp_w*0 +:temp_w] = v339obus[temp_w*0 +:temp_w];
assign v339ibus[data_w*0 +:data_w] = c219obus[data_w*0 +:data_w];
assign c219ibus[temp_w*1 +:temp_w] = v433obus[temp_w*0 +:temp_w];
assign v433ibus[data_w*0 +:data_w] = c219obus[data_w*1 +:data_w];
assign c219ibus[temp_w*2 +:temp_w] = v492obus[temp_w*1 +:temp_w];
assign v492ibus[data_w*1 +:data_w] = c219obus[data_w*2 +:data_w];
assign c219ibus[temp_w*3 +:temp_w] = v732obus[temp_w*1 +:temp_w];
assign v732ibus[data_w*1 +:data_w] = c219obus[data_w*3 +:data_w];
assign c219ibus[temp_w*4 +:temp_w] = v1083obus[temp_w*1 +:temp_w];
assign v1083ibus[data_w*1 +:data_w] = c219obus[data_w*4 +:data_w];
assign c219ibus[temp_w*5 +:temp_w] = v1371obus[temp_w*1 +:temp_w];
assign v1371ibus[data_w*1 +:data_w] = c219obus[data_w*5 +:data_w];
assign c219ibus[temp_w*6 +:temp_w] = v1467obus[temp_w*0 +:temp_w];
assign v1467ibus[data_w*0 +:data_w] = c219obus[data_w*6 +:data_w];
assign c220ibus[temp_w*0 +:temp_w] = v340obus[temp_w*0 +:temp_w];
assign v340ibus[data_w*0 +:data_w] = c220obus[data_w*0 +:data_w];
assign c220ibus[temp_w*1 +:temp_w] = v434obus[temp_w*0 +:temp_w];
assign v434ibus[data_w*0 +:data_w] = c220obus[data_w*1 +:data_w];
assign c220ibus[temp_w*2 +:temp_w] = v493obus[temp_w*1 +:temp_w];
assign v493ibus[data_w*1 +:data_w] = c220obus[data_w*2 +:data_w];
assign c220ibus[temp_w*3 +:temp_w] = v733obus[temp_w*1 +:temp_w];
assign v733ibus[data_w*1 +:data_w] = c220obus[data_w*3 +:data_w];
assign c220ibus[temp_w*4 +:temp_w] = v1084obus[temp_w*1 +:temp_w];
assign v1084ibus[data_w*1 +:data_w] = c220obus[data_w*4 +:data_w];
assign c220ibus[temp_w*5 +:temp_w] = v1372obus[temp_w*1 +:temp_w];
assign v1372ibus[data_w*1 +:data_w] = c220obus[data_w*5 +:data_w];
assign c220ibus[temp_w*6 +:temp_w] = v1468obus[temp_w*0 +:temp_w];
assign v1468ibus[data_w*0 +:data_w] = c220obus[data_w*6 +:data_w];
assign c221ibus[temp_w*0 +:temp_w] = v341obus[temp_w*0 +:temp_w];
assign v341ibus[data_w*0 +:data_w] = c221obus[data_w*0 +:data_w];
assign c221ibus[temp_w*1 +:temp_w] = v435obus[temp_w*0 +:temp_w];
assign v435ibus[data_w*0 +:data_w] = c221obus[data_w*1 +:data_w];
assign c221ibus[temp_w*2 +:temp_w] = v494obus[temp_w*1 +:temp_w];
assign v494ibus[data_w*1 +:data_w] = c221obus[data_w*2 +:data_w];
assign c221ibus[temp_w*3 +:temp_w] = v734obus[temp_w*1 +:temp_w];
assign v734ibus[data_w*1 +:data_w] = c221obus[data_w*3 +:data_w];
assign c221ibus[temp_w*4 +:temp_w] = v1085obus[temp_w*1 +:temp_w];
assign v1085ibus[data_w*1 +:data_w] = c221obus[data_w*4 +:data_w];
assign c221ibus[temp_w*5 +:temp_w] = v1373obus[temp_w*1 +:temp_w];
assign v1373ibus[data_w*1 +:data_w] = c221obus[data_w*5 +:data_w];
assign c221ibus[temp_w*6 +:temp_w] = v1469obus[temp_w*0 +:temp_w];
assign v1469ibus[data_w*0 +:data_w] = c221obus[data_w*6 +:data_w];
assign c222ibus[temp_w*0 +:temp_w] = v342obus[temp_w*0 +:temp_w];
assign v342ibus[data_w*0 +:data_w] = c222obus[data_w*0 +:data_w];
assign c222ibus[temp_w*1 +:temp_w] = v436obus[temp_w*0 +:temp_w];
assign v436ibus[data_w*0 +:data_w] = c222obus[data_w*1 +:data_w];
assign c222ibus[temp_w*2 +:temp_w] = v495obus[temp_w*1 +:temp_w];
assign v495ibus[data_w*1 +:data_w] = c222obus[data_w*2 +:data_w];
assign c222ibus[temp_w*3 +:temp_w] = v735obus[temp_w*1 +:temp_w];
assign v735ibus[data_w*1 +:data_w] = c222obus[data_w*3 +:data_w];
assign c222ibus[temp_w*4 +:temp_w] = v1086obus[temp_w*1 +:temp_w];
assign v1086ibus[data_w*1 +:data_w] = c222obus[data_w*4 +:data_w];
assign c222ibus[temp_w*5 +:temp_w] = v1374obus[temp_w*1 +:temp_w];
assign v1374ibus[data_w*1 +:data_w] = c222obus[data_w*5 +:data_w];
assign c222ibus[temp_w*6 +:temp_w] = v1470obus[temp_w*0 +:temp_w];
assign v1470ibus[data_w*0 +:data_w] = c222obus[data_w*6 +:data_w];
assign c223ibus[temp_w*0 +:temp_w] = v343obus[temp_w*0 +:temp_w];
assign v343ibus[data_w*0 +:data_w] = c223obus[data_w*0 +:data_w];
assign c223ibus[temp_w*1 +:temp_w] = v437obus[temp_w*0 +:temp_w];
assign v437ibus[data_w*0 +:data_w] = c223obus[data_w*1 +:data_w];
assign c223ibus[temp_w*2 +:temp_w] = v496obus[temp_w*1 +:temp_w];
assign v496ibus[data_w*1 +:data_w] = c223obus[data_w*2 +:data_w];
assign c223ibus[temp_w*3 +:temp_w] = v736obus[temp_w*1 +:temp_w];
assign v736ibus[data_w*1 +:data_w] = c223obus[data_w*3 +:data_w];
assign c223ibus[temp_w*4 +:temp_w] = v1087obus[temp_w*1 +:temp_w];
assign v1087ibus[data_w*1 +:data_w] = c223obus[data_w*4 +:data_w];
assign c223ibus[temp_w*5 +:temp_w] = v1375obus[temp_w*1 +:temp_w];
assign v1375ibus[data_w*1 +:data_w] = c223obus[data_w*5 +:data_w];
assign c223ibus[temp_w*6 +:temp_w] = v1471obus[temp_w*0 +:temp_w];
assign v1471ibus[data_w*0 +:data_w] = c223obus[data_w*6 +:data_w];
assign c224ibus[temp_w*0 +:temp_w] = v344obus[temp_w*0 +:temp_w];
assign v344ibus[data_w*0 +:data_w] = c224obus[data_w*0 +:data_w];
assign c224ibus[temp_w*1 +:temp_w] = v438obus[temp_w*0 +:temp_w];
assign v438ibus[data_w*0 +:data_w] = c224obus[data_w*1 +:data_w];
assign c224ibus[temp_w*2 +:temp_w] = v497obus[temp_w*1 +:temp_w];
assign v497ibus[data_w*1 +:data_w] = c224obus[data_w*2 +:data_w];
assign c224ibus[temp_w*3 +:temp_w] = v737obus[temp_w*1 +:temp_w];
assign v737ibus[data_w*1 +:data_w] = c224obus[data_w*3 +:data_w];
assign c224ibus[temp_w*4 +:temp_w] = v1088obus[temp_w*1 +:temp_w];
assign v1088ibus[data_w*1 +:data_w] = c224obus[data_w*4 +:data_w];
assign c224ibus[temp_w*5 +:temp_w] = v1376obus[temp_w*1 +:temp_w];
assign v1376ibus[data_w*1 +:data_w] = c224obus[data_w*5 +:data_w];
assign c224ibus[temp_w*6 +:temp_w] = v1472obus[temp_w*0 +:temp_w];
assign v1472ibus[data_w*0 +:data_w] = c224obus[data_w*6 +:data_w];
assign c225ibus[temp_w*0 +:temp_w] = v345obus[temp_w*0 +:temp_w];
assign v345ibus[data_w*0 +:data_w] = c225obus[data_w*0 +:data_w];
assign c225ibus[temp_w*1 +:temp_w] = v439obus[temp_w*0 +:temp_w];
assign v439ibus[data_w*0 +:data_w] = c225obus[data_w*1 +:data_w];
assign c225ibus[temp_w*2 +:temp_w] = v498obus[temp_w*1 +:temp_w];
assign v498ibus[data_w*1 +:data_w] = c225obus[data_w*2 +:data_w];
assign c225ibus[temp_w*3 +:temp_w] = v738obus[temp_w*1 +:temp_w];
assign v738ibus[data_w*1 +:data_w] = c225obus[data_w*3 +:data_w];
assign c225ibus[temp_w*4 +:temp_w] = v1089obus[temp_w*1 +:temp_w];
assign v1089ibus[data_w*1 +:data_w] = c225obus[data_w*4 +:data_w];
assign c225ibus[temp_w*5 +:temp_w] = v1377obus[temp_w*1 +:temp_w];
assign v1377ibus[data_w*1 +:data_w] = c225obus[data_w*5 +:data_w];
assign c225ibus[temp_w*6 +:temp_w] = v1473obus[temp_w*0 +:temp_w];
assign v1473ibus[data_w*0 +:data_w] = c225obus[data_w*6 +:data_w];
assign c226ibus[temp_w*0 +:temp_w] = v346obus[temp_w*0 +:temp_w];
assign v346ibus[data_w*0 +:data_w] = c226obus[data_w*0 +:data_w];
assign c226ibus[temp_w*1 +:temp_w] = v440obus[temp_w*0 +:temp_w];
assign v440ibus[data_w*0 +:data_w] = c226obus[data_w*1 +:data_w];
assign c226ibus[temp_w*2 +:temp_w] = v499obus[temp_w*1 +:temp_w];
assign v499ibus[data_w*1 +:data_w] = c226obus[data_w*2 +:data_w];
assign c226ibus[temp_w*3 +:temp_w] = v739obus[temp_w*1 +:temp_w];
assign v739ibus[data_w*1 +:data_w] = c226obus[data_w*3 +:data_w];
assign c226ibus[temp_w*4 +:temp_w] = v1090obus[temp_w*1 +:temp_w];
assign v1090ibus[data_w*1 +:data_w] = c226obus[data_w*4 +:data_w];
assign c226ibus[temp_w*5 +:temp_w] = v1378obus[temp_w*1 +:temp_w];
assign v1378ibus[data_w*1 +:data_w] = c226obus[data_w*5 +:data_w];
assign c226ibus[temp_w*6 +:temp_w] = v1474obus[temp_w*0 +:temp_w];
assign v1474ibus[data_w*0 +:data_w] = c226obus[data_w*6 +:data_w];
assign c227ibus[temp_w*0 +:temp_w] = v347obus[temp_w*0 +:temp_w];
assign v347ibus[data_w*0 +:data_w] = c227obus[data_w*0 +:data_w];
assign c227ibus[temp_w*1 +:temp_w] = v441obus[temp_w*0 +:temp_w];
assign v441ibus[data_w*0 +:data_w] = c227obus[data_w*1 +:data_w];
assign c227ibus[temp_w*2 +:temp_w] = v500obus[temp_w*1 +:temp_w];
assign v500ibus[data_w*1 +:data_w] = c227obus[data_w*2 +:data_w];
assign c227ibus[temp_w*3 +:temp_w] = v740obus[temp_w*1 +:temp_w];
assign v740ibus[data_w*1 +:data_w] = c227obus[data_w*3 +:data_w];
assign c227ibus[temp_w*4 +:temp_w] = v1091obus[temp_w*1 +:temp_w];
assign v1091ibus[data_w*1 +:data_w] = c227obus[data_w*4 +:data_w];
assign c227ibus[temp_w*5 +:temp_w] = v1379obus[temp_w*1 +:temp_w];
assign v1379ibus[data_w*1 +:data_w] = c227obus[data_w*5 +:data_w];
assign c227ibus[temp_w*6 +:temp_w] = v1475obus[temp_w*0 +:temp_w];
assign v1475ibus[data_w*0 +:data_w] = c227obus[data_w*6 +:data_w];
assign c228ibus[temp_w*0 +:temp_w] = v348obus[temp_w*0 +:temp_w];
assign v348ibus[data_w*0 +:data_w] = c228obus[data_w*0 +:data_w];
assign c228ibus[temp_w*1 +:temp_w] = v442obus[temp_w*0 +:temp_w];
assign v442ibus[data_w*0 +:data_w] = c228obus[data_w*1 +:data_w];
assign c228ibus[temp_w*2 +:temp_w] = v501obus[temp_w*1 +:temp_w];
assign v501ibus[data_w*1 +:data_w] = c228obus[data_w*2 +:data_w];
assign c228ibus[temp_w*3 +:temp_w] = v741obus[temp_w*1 +:temp_w];
assign v741ibus[data_w*1 +:data_w] = c228obus[data_w*3 +:data_w];
assign c228ibus[temp_w*4 +:temp_w] = v1092obus[temp_w*1 +:temp_w];
assign v1092ibus[data_w*1 +:data_w] = c228obus[data_w*4 +:data_w];
assign c228ibus[temp_w*5 +:temp_w] = v1380obus[temp_w*1 +:temp_w];
assign v1380ibus[data_w*1 +:data_w] = c228obus[data_w*5 +:data_w];
assign c228ibus[temp_w*6 +:temp_w] = v1476obus[temp_w*0 +:temp_w];
assign v1476ibus[data_w*0 +:data_w] = c228obus[data_w*6 +:data_w];
assign c229ibus[temp_w*0 +:temp_w] = v349obus[temp_w*0 +:temp_w];
assign v349ibus[data_w*0 +:data_w] = c229obus[data_w*0 +:data_w];
assign c229ibus[temp_w*1 +:temp_w] = v443obus[temp_w*0 +:temp_w];
assign v443ibus[data_w*0 +:data_w] = c229obus[data_w*1 +:data_w];
assign c229ibus[temp_w*2 +:temp_w] = v502obus[temp_w*1 +:temp_w];
assign v502ibus[data_w*1 +:data_w] = c229obus[data_w*2 +:data_w];
assign c229ibus[temp_w*3 +:temp_w] = v742obus[temp_w*1 +:temp_w];
assign v742ibus[data_w*1 +:data_w] = c229obus[data_w*3 +:data_w];
assign c229ibus[temp_w*4 +:temp_w] = v1093obus[temp_w*1 +:temp_w];
assign v1093ibus[data_w*1 +:data_w] = c229obus[data_w*4 +:data_w];
assign c229ibus[temp_w*5 +:temp_w] = v1381obus[temp_w*1 +:temp_w];
assign v1381ibus[data_w*1 +:data_w] = c229obus[data_w*5 +:data_w];
assign c229ibus[temp_w*6 +:temp_w] = v1477obus[temp_w*0 +:temp_w];
assign v1477ibus[data_w*0 +:data_w] = c229obus[data_w*6 +:data_w];
assign c230ibus[temp_w*0 +:temp_w] = v350obus[temp_w*0 +:temp_w];
assign v350ibus[data_w*0 +:data_w] = c230obus[data_w*0 +:data_w];
assign c230ibus[temp_w*1 +:temp_w] = v444obus[temp_w*0 +:temp_w];
assign v444ibus[data_w*0 +:data_w] = c230obus[data_w*1 +:data_w];
assign c230ibus[temp_w*2 +:temp_w] = v503obus[temp_w*1 +:temp_w];
assign v503ibus[data_w*1 +:data_w] = c230obus[data_w*2 +:data_w];
assign c230ibus[temp_w*3 +:temp_w] = v743obus[temp_w*1 +:temp_w];
assign v743ibus[data_w*1 +:data_w] = c230obus[data_w*3 +:data_w];
assign c230ibus[temp_w*4 +:temp_w] = v1094obus[temp_w*1 +:temp_w];
assign v1094ibus[data_w*1 +:data_w] = c230obus[data_w*4 +:data_w];
assign c230ibus[temp_w*5 +:temp_w] = v1382obus[temp_w*1 +:temp_w];
assign v1382ibus[data_w*1 +:data_w] = c230obus[data_w*5 +:data_w];
assign c230ibus[temp_w*6 +:temp_w] = v1478obus[temp_w*0 +:temp_w];
assign v1478ibus[data_w*0 +:data_w] = c230obus[data_w*6 +:data_w];
assign c231ibus[temp_w*0 +:temp_w] = v351obus[temp_w*0 +:temp_w];
assign v351ibus[data_w*0 +:data_w] = c231obus[data_w*0 +:data_w];
assign c231ibus[temp_w*1 +:temp_w] = v445obus[temp_w*0 +:temp_w];
assign v445ibus[data_w*0 +:data_w] = c231obus[data_w*1 +:data_w];
assign c231ibus[temp_w*2 +:temp_w] = v504obus[temp_w*1 +:temp_w];
assign v504ibus[data_w*1 +:data_w] = c231obus[data_w*2 +:data_w];
assign c231ibus[temp_w*3 +:temp_w] = v744obus[temp_w*1 +:temp_w];
assign v744ibus[data_w*1 +:data_w] = c231obus[data_w*3 +:data_w];
assign c231ibus[temp_w*4 +:temp_w] = v1095obus[temp_w*1 +:temp_w];
assign v1095ibus[data_w*1 +:data_w] = c231obus[data_w*4 +:data_w];
assign c231ibus[temp_w*5 +:temp_w] = v1383obus[temp_w*1 +:temp_w];
assign v1383ibus[data_w*1 +:data_w] = c231obus[data_w*5 +:data_w];
assign c231ibus[temp_w*6 +:temp_w] = v1479obus[temp_w*0 +:temp_w];
assign v1479ibus[data_w*0 +:data_w] = c231obus[data_w*6 +:data_w];
assign c232ibus[temp_w*0 +:temp_w] = v352obus[temp_w*0 +:temp_w];
assign v352ibus[data_w*0 +:data_w] = c232obus[data_w*0 +:data_w];
assign c232ibus[temp_w*1 +:temp_w] = v446obus[temp_w*0 +:temp_w];
assign v446ibus[data_w*0 +:data_w] = c232obus[data_w*1 +:data_w];
assign c232ibus[temp_w*2 +:temp_w] = v505obus[temp_w*1 +:temp_w];
assign v505ibus[data_w*1 +:data_w] = c232obus[data_w*2 +:data_w];
assign c232ibus[temp_w*3 +:temp_w] = v745obus[temp_w*1 +:temp_w];
assign v745ibus[data_w*1 +:data_w] = c232obus[data_w*3 +:data_w];
assign c232ibus[temp_w*4 +:temp_w] = v1096obus[temp_w*1 +:temp_w];
assign v1096ibus[data_w*1 +:data_w] = c232obus[data_w*4 +:data_w];
assign c232ibus[temp_w*5 +:temp_w] = v1384obus[temp_w*1 +:temp_w];
assign v1384ibus[data_w*1 +:data_w] = c232obus[data_w*5 +:data_w];
assign c232ibus[temp_w*6 +:temp_w] = v1480obus[temp_w*0 +:temp_w];
assign v1480ibus[data_w*0 +:data_w] = c232obus[data_w*6 +:data_w];
assign c233ibus[temp_w*0 +:temp_w] = v353obus[temp_w*0 +:temp_w];
assign v353ibus[data_w*0 +:data_w] = c233obus[data_w*0 +:data_w];
assign c233ibus[temp_w*1 +:temp_w] = v447obus[temp_w*0 +:temp_w];
assign v447ibus[data_w*0 +:data_w] = c233obus[data_w*1 +:data_w];
assign c233ibus[temp_w*2 +:temp_w] = v506obus[temp_w*1 +:temp_w];
assign v506ibus[data_w*1 +:data_w] = c233obus[data_w*2 +:data_w];
assign c233ibus[temp_w*3 +:temp_w] = v746obus[temp_w*1 +:temp_w];
assign v746ibus[data_w*1 +:data_w] = c233obus[data_w*3 +:data_w];
assign c233ibus[temp_w*4 +:temp_w] = v1097obus[temp_w*1 +:temp_w];
assign v1097ibus[data_w*1 +:data_w] = c233obus[data_w*4 +:data_w];
assign c233ibus[temp_w*5 +:temp_w] = v1385obus[temp_w*1 +:temp_w];
assign v1385ibus[data_w*1 +:data_w] = c233obus[data_w*5 +:data_w];
assign c233ibus[temp_w*6 +:temp_w] = v1481obus[temp_w*0 +:temp_w];
assign v1481ibus[data_w*0 +:data_w] = c233obus[data_w*6 +:data_w];
assign c234ibus[temp_w*0 +:temp_w] = v354obus[temp_w*0 +:temp_w];
assign v354ibus[data_w*0 +:data_w] = c234obus[data_w*0 +:data_w];
assign c234ibus[temp_w*1 +:temp_w] = v448obus[temp_w*0 +:temp_w];
assign v448ibus[data_w*0 +:data_w] = c234obus[data_w*1 +:data_w];
assign c234ibus[temp_w*2 +:temp_w] = v507obus[temp_w*1 +:temp_w];
assign v507ibus[data_w*1 +:data_w] = c234obus[data_w*2 +:data_w];
assign c234ibus[temp_w*3 +:temp_w] = v747obus[temp_w*1 +:temp_w];
assign v747ibus[data_w*1 +:data_w] = c234obus[data_w*3 +:data_w];
assign c234ibus[temp_w*4 +:temp_w] = v1098obus[temp_w*1 +:temp_w];
assign v1098ibus[data_w*1 +:data_w] = c234obus[data_w*4 +:data_w];
assign c234ibus[temp_w*5 +:temp_w] = v1386obus[temp_w*1 +:temp_w];
assign v1386ibus[data_w*1 +:data_w] = c234obus[data_w*5 +:data_w];
assign c234ibus[temp_w*6 +:temp_w] = v1482obus[temp_w*0 +:temp_w];
assign v1482ibus[data_w*0 +:data_w] = c234obus[data_w*6 +:data_w];
assign c235ibus[temp_w*0 +:temp_w] = v355obus[temp_w*0 +:temp_w];
assign v355ibus[data_w*0 +:data_w] = c235obus[data_w*0 +:data_w];
assign c235ibus[temp_w*1 +:temp_w] = v449obus[temp_w*0 +:temp_w];
assign v449ibus[data_w*0 +:data_w] = c235obus[data_w*1 +:data_w];
assign c235ibus[temp_w*2 +:temp_w] = v508obus[temp_w*1 +:temp_w];
assign v508ibus[data_w*1 +:data_w] = c235obus[data_w*2 +:data_w];
assign c235ibus[temp_w*3 +:temp_w] = v748obus[temp_w*1 +:temp_w];
assign v748ibus[data_w*1 +:data_w] = c235obus[data_w*3 +:data_w];
assign c235ibus[temp_w*4 +:temp_w] = v1099obus[temp_w*1 +:temp_w];
assign v1099ibus[data_w*1 +:data_w] = c235obus[data_w*4 +:data_w];
assign c235ibus[temp_w*5 +:temp_w] = v1387obus[temp_w*1 +:temp_w];
assign v1387ibus[data_w*1 +:data_w] = c235obus[data_w*5 +:data_w];
assign c235ibus[temp_w*6 +:temp_w] = v1483obus[temp_w*0 +:temp_w];
assign v1483ibus[data_w*0 +:data_w] = c235obus[data_w*6 +:data_w];
assign c236ibus[temp_w*0 +:temp_w] = v356obus[temp_w*0 +:temp_w];
assign v356ibus[data_w*0 +:data_w] = c236obus[data_w*0 +:data_w];
assign c236ibus[temp_w*1 +:temp_w] = v450obus[temp_w*0 +:temp_w];
assign v450ibus[data_w*0 +:data_w] = c236obus[data_w*1 +:data_w];
assign c236ibus[temp_w*2 +:temp_w] = v509obus[temp_w*1 +:temp_w];
assign v509ibus[data_w*1 +:data_w] = c236obus[data_w*2 +:data_w];
assign c236ibus[temp_w*3 +:temp_w] = v749obus[temp_w*1 +:temp_w];
assign v749ibus[data_w*1 +:data_w] = c236obus[data_w*3 +:data_w];
assign c236ibus[temp_w*4 +:temp_w] = v1100obus[temp_w*1 +:temp_w];
assign v1100ibus[data_w*1 +:data_w] = c236obus[data_w*4 +:data_w];
assign c236ibus[temp_w*5 +:temp_w] = v1388obus[temp_w*1 +:temp_w];
assign v1388ibus[data_w*1 +:data_w] = c236obus[data_w*5 +:data_w];
assign c236ibus[temp_w*6 +:temp_w] = v1484obus[temp_w*0 +:temp_w];
assign v1484ibus[data_w*0 +:data_w] = c236obus[data_w*6 +:data_w];
assign c237ibus[temp_w*0 +:temp_w] = v357obus[temp_w*0 +:temp_w];
assign v357ibus[data_w*0 +:data_w] = c237obus[data_w*0 +:data_w];
assign c237ibus[temp_w*1 +:temp_w] = v451obus[temp_w*0 +:temp_w];
assign v451ibus[data_w*0 +:data_w] = c237obus[data_w*1 +:data_w];
assign c237ibus[temp_w*2 +:temp_w] = v510obus[temp_w*1 +:temp_w];
assign v510ibus[data_w*1 +:data_w] = c237obus[data_w*2 +:data_w];
assign c237ibus[temp_w*3 +:temp_w] = v750obus[temp_w*1 +:temp_w];
assign v750ibus[data_w*1 +:data_w] = c237obus[data_w*3 +:data_w];
assign c237ibus[temp_w*4 +:temp_w] = v1101obus[temp_w*1 +:temp_w];
assign v1101ibus[data_w*1 +:data_w] = c237obus[data_w*4 +:data_w];
assign c237ibus[temp_w*5 +:temp_w] = v1389obus[temp_w*1 +:temp_w];
assign v1389ibus[data_w*1 +:data_w] = c237obus[data_w*5 +:data_w];
assign c237ibus[temp_w*6 +:temp_w] = v1485obus[temp_w*0 +:temp_w];
assign v1485ibus[data_w*0 +:data_w] = c237obus[data_w*6 +:data_w];
assign c238ibus[temp_w*0 +:temp_w] = v358obus[temp_w*0 +:temp_w];
assign v358ibus[data_w*0 +:data_w] = c238obus[data_w*0 +:data_w];
assign c238ibus[temp_w*1 +:temp_w] = v452obus[temp_w*0 +:temp_w];
assign v452ibus[data_w*0 +:data_w] = c238obus[data_w*1 +:data_w];
assign c238ibus[temp_w*2 +:temp_w] = v511obus[temp_w*1 +:temp_w];
assign v511ibus[data_w*1 +:data_w] = c238obus[data_w*2 +:data_w];
assign c238ibus[temp_w*3 +:temp_w] = v751obus[temp_w*1 +:temp_w];
assign v751ibus[data_w*1 +:data_w] = c238obus[data_w*3 +:data_w];
assign c238ibus[temp_w*4 +:temp_w] = v1102obus[temp_w*1 +:temp_w];
assign v1102ibus[data_w*1 +:data_w] = c238obus[data_w*4 +:data_w];
assign c238ibus[temp_w*5 +:temp_w] = v1390obus[temp_w*1 +:temp_w];
assign v1390ibus[data_w*1 +:data_w] = c238obus[data_w*5 +:data_w];
assign c238ibus[temp_w*6 +:temp_w] = v1486obus[temp_w*0 +:temp_w];
assign v1486ibus[data_w*0 +:data_w] = c238obus[data_w*6 +:data_w];
assign c239ibus[temp_w*0 +:temp_w] = v359obus[temp_w*0 +:temp_w];
assign v359ibus[data_w*0 +:data_w] = c239obus[data_w*0 +:data_w];
assign c239ibus[temp_w*1 +:temp_w] = v453obus[temp_w*0 +:temp_w];
assign v453ibus[data_w*0 +:data_w] = c239obus[data_w*1 +:data_w];
assign c239ibus[temp_w*2 +:temp_w] = v512obus[temp_w*1 +:temp_w];
assign v512ibus[data_w*1 +:data_w] = c239obus[data_w*2 +:data_w];
assign c239ibus[temp_w*3 +:temp_w] = v752obus[temp_w*1 +:temp_w];
assign v752ibus[data_w*1 +:data_w] = c239obus[data_w*3 +:data_w];
assign c239ibus[temp_w*4 +:temp_w] = v1103obus[temp_w*1 +:temp_w];
assign v1103ibus[data_w*1 +:data_w] = c239obus[data_w*4 +:data_w];
assign c239ibus[temp_w*5 +:temp_w] = v1391obus[temp_w*1 +:temp_w];
assign v1391ibus[data_w*1 +:data_w] = c239obus[data_w*5 +:data_w];
assign c239ibus[temp_w*6 +:temp_w] = v1487obus[temp_w*0 +:temp_w];
assign v1487ibus[data_w*0 +:data_w] = c239obus[data_w*6 +:data_w];
assign c240ibus[temp_w*0 +:temp_w] = v360obus[temp_w*0 +:temp_w];
assign v360ibus[data_w*0 +:data_w] = c240obus[data_w*0 +:data_w];
assign c240ibus[temp_w*1 +:temp_w] = v454obus[temp_w*0 +:temp_w];
assign v454ibus[data_w*0 +:data_w] = c240obus[data_w*1 +:data_w];
assign c240ibus[temp_w*2 +:temp_w] = v513obus[temp_w*1 +:temp_w];
assign v513ibus[data_w*1 +:data_w] = c240obus[data_w*2 +:data_w];
assign c240ibus[temp_w*3 +:temp_w] = v753obus[temp_w*1 +:temp_w];
assign v753ibus[data_w*1 +:data_w] = c240obus[data_w*3 +:data_w];
assign c240ibus[temp_w*4 +:temp_w] = v1104obus[temp_w*1 +:temp_w];
assign v1104ibus[data_w*1 +:data_w] = c240obus[data_w*4 +:data_w];
assign c240ibus[temp_w*5 +:temp_w] = v1392obus[temp_w*1 +:temp_w];
assign v1392ibus[data_w*1 +:data_w] = c240obus[data_w*5 +:data_w];
assign c240ibus[temp_w*6 +:temp_w] = v1488obus[temp_w*0 +:temp_w];
assign v1488ibus[data_w*0 +:data_w] = c240obus[data_w*6 +:data_w];
assign c241ibus[temp_w*0 +:temp_w] = v361obus[temp_w*0 +:temp_w];
assign v361ibus[data_w*0 +:data_w] = c241obus[data_w*0 +:data_w];
assign c241ibus[temp_w*1 +:temp_w] = v455obus[temp_w*0 +:temp_w];
assign v455ibus[data_w*0 +:data_w] = c241obus[data_w*1 +:data_w];
assign c241ibus[temp_w*2 +:temp_w] = v514obus[temp_w*1 +:temp_w];
assign v514ibus[data_w*1 +:data_w] = c241obus[data_w*2 +:data_w];
assign c241ibus[temp_w*3 +:temp_w] = v754obus[temp_w*1 +:temp_w];
assign v754ibus[data_w*1 +:data_w] = c241obus[data_w*3 +:data_w];
assign c241ibus[temp_w*4 +:temp_w] = v1105obus[temp_w*1 +:temp_w];
assign v1105ibus[data_w*1 +:data_w] = c241obus[data_w*4 +:data_w];
assign c241ibus[temp_w*5 +:temp_w] = v1393obus[temp_w*1 +:temp_w];
assign v1393ibus[data_w*1 +:data_w] = c241obus[data_w*5 +:data_w];
assign c241ibus[temp_w*6 +:temp_w] = v1489obus[temp_w*0 +:temp_w];
assign v1489ibus[data_w*0 +:data_w] = c241obus[data_w*6 +:data_w];
assign c242ibus[temp_w*0 +:temp_w] = v362obus[temp_w*0 +:temp_w];
assign v362ibus[data_w*0 +:data_w] = c242obus[data_w*0 +:data_w];
assign c242ibus[temp_w*1 +:temp_w] = v456obus[temp_w*0 +:temp_w];
assign v456ibus[data_w*0 +:data_w] = c242obus[data_w*1 +:data_w];
assign c242ibus[temp_w*2 +:temp_w] = v515obus[temp_w*1 +:temp_w];
assign v515ibus[data_w*1 +:data_w] = c242obus[data_w*2 +:data_w];
assign c242ibus[temp_w*3 +:temp_w] = v755obus[temp_w*1 +:temp_w];
assign v755ibus[data_w*1 +:data_w] = c242obus[data_w*3 +:data_w];
assign c242ibus[temp_w*4 +:temp_w] = v1106obus[temp_w*1 +:temp_w];
assign v1106ibus[data_w*1 +:data_w] = c242obus[data_w*4 +:data_w];
assign c242ibus[temp_w*5 +:temp_w] = v1394obus[temp_w*1 +:temp_w];
assign v1394ibus[data_w*1 +:data_w] = c242obus[data_w*5 +:data_w];
assign c242ibus[temp_w*6 +:temp_w] = v1490obus[temp_w*0 +:temp_w];
assign v1490ibus[data_w*0 +:data_w] = c242obus[data_w*6 +:data_w];
assign c243ibus[temp_w*0 +:temp_w] = v363obus[temp_w*0 +:temp_w];
assign v363ibus[data_w*0 +:data_w] = c243obus[data_w*0 +:data_w];
assign c243ibus[temp_w*1 +:temp_w] = v457obus[temp_w*0 +:temp_w];
assign v457ibus[data_w*0 +:data_w] = c243obus[data_w*1 +:data_w];
assign c243ibus[temp_w*2 +:temp_w] = v516obus[temp_w*1 +:temp_w];
assign v516ibus[data_w*1 +:data_w] = c243obus[data_w*2 +:data_w];
assign c243ibus[temp_w*3 +:temp_w] = v756obus[temp_w*1 +:temp_w];
assign v756ibus[data_w*1 +:data_w] = c243obus[data_w*3 +:data_w];
assign c243ibus[temp_w*4 +:temp_w] = v1107obus[temp_w*1 +:temp_w];
assign v1107ibus[data_w*1 +:data_w] = c243obus[data_w*4 +:data_w];
assign c243ibus[temp_w*5 +:temp_w] = v1395obus[temp_w*1 +:temp_w];
assign v1395ibus[data_w*1 +:data_w] = c243obus[data_w*5 +:data_w];
assign c243ibus[temp_w*6 +:temp_w] = v1491obus[temp_w*0 +:temp_w];
assign v1491ibus[data_w*0 +:data_w] = c243obus[data_w*6 +:data_w];
assign c244ibus[temp_w*0 +:temp_w] = v364obus[temp_w*0 +:temp_w];
assign v364ibus[data_w*0 +:data_w] = c244obus[data_w*0 +:data_w];
assign c244ibus[temp_w*1 +:temp_w] = v458obus[temp_w*0 +:temp_w];
assign v458ibus[data_w*0 +:data_w] = c244obus[data_w*1 +:data_w];
assign c244ibus[temp_w*2 +:temp_w] = v517obus[temp_w*1 +:temp_w];
assign v517ibus[data_w*1 +:data_w] = c244obus[data_w*2 +:data_w];
assign c244ibus[temp_w*3 +:temp_w] = v757obus[temp_w*1 +:temp_w];
assign v757ibus[data_w*1 +:data_w] = c244obus[data_w*3 +:data_w];
assign c244ibus[temp_w*4 +:temp_w] = v1108obus[temp_w*1 +:temp_w];
assign v1108ibus[data_w*1 +:data_w] = c244obus[data_w*4 +:data_w];
assign c244ibus[temp_w*5 +:temp_w] = v1396obus[temp_w*1 +:temp_w];
assign v1396ibus[data_w*1 +:data_w] = c244obus[data_w*5 +:data_w];
assign c244ibus[temp_w*6 +:temp_w] = v1492obus[temp_w*0 +:temp_w];
assign v1492ibus[data_w*0 +:data_w] = c244obus[data_w*6 +:data_w];
assign c245ibus[temp_w*0 +:temp_w] = v365obus[temp_w*0 +:temp_w];
assign v365ibus[data_w*0 +:data_w] = c245obus[data_w*0 +:data_w];
assign c245ibus[temp_w*1 +:temp_w] = v459obus[temp_w*0 +:temp_w];
assign v459ibus[data_w*0 +:data_w] = c245obus[data_w*1 +:data_w];
assign c245ibus[temp_w*2 +:temp_w] = v518obus[temp_w*1 +:temp_w];
assign v518ibus[data_w*1 +:data_w] = c245obus[data_w*2 +:data_w];
assign c245ibus[temp_w*3 +:temp_w] = v758obus[temp_w*1 +:temp_w];
assign v758ibus[data_w*1 +:data_w] = c245obus[data_w*3 +:data_w];
assign c245ibus[temp_w*4 +:temp_w] = v1109obus[temp_w*1 +:temp_w];
assign v1109ibus[data_w*1 +:data_w] = c245obus[data_w*4 +:data_w];
assign c245ibus[temp_w*5 +:temp_w] = v1397obus[temp_w*1 +:temp_w];
assign v1397ibus[data_w*1 +:data_w] = c245obus[data_w*5 +:data_w];
assign c245ibus[temp_w*6 +:temp_w] = v1493obus[temp_w*0 +:temp_w];
assign v1493ibus[data_w*0 +:data_w] = c245obus[data_w*6 +:data_w];
assign c246ibus[temp_w*0 +:temp_w] = v366obus[temp_w*0 +:temp_w];
assign v366ibus[data_w*0 +:data_w] = c246obus[data_w*0 +:data_w];
assign c246ibus[temp_w*1 +:temp_w] = v460obus[temp_w*0 +:temp_w];
assign v460ibus[data_w*0 +:data_w] = c246obus[data_w*1 +:data_w];
assign c246ibus[temp_w*2 +:temp_w] = v519obus[temp_w*1 +:temp_w];
assign v519ibus[data_w*1 +:data_w] = c246obus[data_w*2 +:data_w];
assign c246ibus[temp_w*3 +:temp_w] = v759obus[temp_w*1 +:temp_w];
assign v759ibus[data_w*1 +:data_w] = c246obus[data_w*3 +:data_w];
assign c246ibus[temp_w*4 +:temp_w] = v1110obus[temp_w*1 +:temp_w];
assign v1110ibus[data_w*1 +:data_w] = c246obus[data_w*4 +:data_w];
assign c246ibus[temp_w*5 +:temp_w] = v1398obus[temp_w*1 +:temp_w];
assign v1398ibus[data_w*1 +:data_w] = c246obus[data_w*5 +:data_w];
assign c246ibus[temp_w*6 +:temp_w] = v1494obus[temp_w*0 +:temp_w];
assign v1494ibus[data_w*0 +:data_w] = c246obus[data_w*6 +:data_w];
assign c247ibus[temp_w*0 +:temp_w] = v367obus[temp_w*0 +:temp_w];
assign v367ibus[data_w*0 +:data_w] = c247obus[data_w*0 +:data_w];
assign c247ibus[temp_w*1 +:temp_w] = v461obus[temp_w*0 +:temp_w];
assign v461ibus[data_w*0 +:data_w] = c247obus[data_w*1 +:data_w];
assign c247ibus[temp_w*2 +:temp_w] = v520obus[temp_w*1 +:temp_w];
assign v520ibus[data_w*1 +:data_w] = c247obus[data_w*2 +:data_w];
assign c247ibus[temp_w*3 +:temp_w] = v760obus[temp_w*1 +:temp_w];
assign v760ibus[data_w*1 +:data_w] = c247obus[data_w*3 +:data_w];
assign c247ibus[temp_w*4 +:temp_w] = v1111obus[temp_w*1 +:temp_w];
assign v1111ibus[data_w*1 +:data_w] = c247obus[data_w*4 +:data_w];
assign c247ibus[temp_w*5 +:temp_w] = v1399obus[temp_w*1 +:temp_w];
assign v1399ibus[data_w*1 +:data_w] = c247obus[data_w*5 +:data_w];
assign c247ibus[temp_w*6 +:temp_w] = v1495obus[temp_w*0 +:temp_w];
assign v1495ibus[data_w*0 +:data_w] = c247obus[data_w*6 +:data_w];
assign c248ibus[temp_w*0 +:temp_w] = v368obus[temp_w*0 +:temp_w];
assign v368ibus[data_w*0 +:data_w] = c248obus[data_w*0 +:data_w];
assign c248ibus[temp_w*1 +:temp_w] = v462obus[temp_w*0 +:temp_w];
assign v462ibus[data_w*0 +:data_w] = c248obus[data_w*1 +:data_w];
assign c248ibus[temp_w*2 +:temp_w] = v521obus[temp_w*1 +:temp_w];
assign v521ibus[data_w*1 +:data_w] = c248obus[data_w*2 +:data_w];
assign c248ibus[temp_w*3 +:temp_w] = v761obus[temp_w*1 +:temp_w];
assign v761ibus[data_w*1 +:data_w] = c248obus[data_w*3 +:data_w];
assign c248ibus[temp_w*4 +:temp_w] = v1112obus[temp_w*1 +:temp_w];
assign v1112ibus[data_w*1 +:data_w] = c248obus[data_w*4 +:data_w];
assign c248ibus[temp_w*5 +:temp_w] = v1400obus[temp_w*1 +:temp_w];
assign v1400ibus[data_w*1 +:data_w] = c248obus[data_w*5 +:data_w];
assign c248ibus[temp_w*6 +:temp_w] = v1496obus[temp_w*0 +:temp_w];
assign v1496ibus[data_w*0 +:data_w] = c248obus[data_w*6 +:data_w];
assign c249ibus[temp_w*0 +:temp_w] = v369obus[temp_w*0 +:temp_w];
assign v369ibus[data_w*0 +:data_w] = c249obus[data_w*0 +:data_w];
assign c249ibus[temp_w*1 +:temp_w] = v463obus[temp_w*0 +:temp_w];
assign v463ibus[data_w*0 +:data_w] = c249obus[data_w*1 +:data_w];
assign c249ibus[temp_w*2 +:temp_w] = v522obus[temp_w*1 +:temp_w];
assign v522ibus[data_w*1 +:data_w] = c249obus[data_w*2 +:data_w];
assign c249ibus[temp_w*3 +:temp_w] = v762obus[temp_w*1 +:temp_w];
assign v762ibus[data_w*1 +:data_w] = c249obus[data_w*3 +:data_w];
assign c249ibus[temp_w*4 +:temp_w] = v1113obus[temp_w*1 +:temp_w];
assign v1113ibus[data_w*1 +:data_w] = c249obus[data_w*4 +:data_w];
assign c249ibus[temp_w*5 +:temp_w] = v1401obus[temp_w*1 +:temp_w];
assign v1401ibus[data_w*1 +:data_w] = c249obus[data_w*5 +:data_w];
assign c249ibus[temp_w*6 +:temp_w] = v1497obus[temp_w*0 +:temp_w];
assign v1497ibus[data_w*0 +:data_w] = c249obus[data_w*6 +:data_w];
assign c250ibus[temp_w*0 +:temp_w] = v370obus[temp_w*0 +:temp_w];
assign v370ibus[data_w*0 +:data_w] = c250obus[data_w*0 +:data_w];
assign c250ibus[temp_w*1 +:temp_w] = v464obus[temp_w*0 +:temp_w];
assign v464ibus[data_w*0 +:data_w] = c250obus[data_w*1 +:data_w];
assign c250ibus[temp_w*2 +:temp_w] = v523obus[temp_w*1 +:temp_w];
assign v523ibus[data_w*1 +:data_w] = c250obus[data_w*2 +:data_w];
assign c250ibus[temp_w*3 +:temp_w] = v763obus[temp_w*1 +:temp_w];
assign v763ibus[data_w*1 +:data_w] = c250obus[data_w*3 +:data_w];
assign c250ibus[temp_w*4 +:temp_w] = v1114obus[temp_w*1 +:temp_w];
assign v1114ibus[data_w*1 +:data_w] = c250obus[data_w*4 +:data_w];
assign c250ibus[temp_w*5 +:temp_w] = v1402obus[temp_w*1 +:temp_w];
assign v1402ibus[data_w*1 +:data_w] = c250obus[data_w*5 +:data_w];
assign c250ibus[temp_w*6 +:temp_w] = v1498obus[temp_w*0 +:temp_w];
assign v1498ibus[data_w*0 +:data_w] = c250obus[data_w*6 +:data_w];
assign c251ibus[temp_w*0 +:temp_w] = v371obus[temp_w*0 +:temp_w];
assign v371ibus[data_w*0 +:data_w] = c251obus[data_w*0 +:data_w];
assign c251ibus[temp_w*1 +:temp_w] = v465obus[temp_w*0 +:temp_w];
assign v465ibus[data_w*0 +:data_w] = c251obus[data_w*1 +:data_w];
assign c251ibus[temp_w*2 +:temp_w] = v524obus[temp_w*1 +:temp_w];
assign v524ibus[data_w*1 +:data_w] = c251obus[data_w*2 +:data_w];
assign c251ibus[temp_w*3 +:temp_w] = v764obus[temp_w*1 +:temp_w];
assign v764ibus[data_w*1 +:data_w] = c251obus[data_w*3 +:data_w];
assign c251ibus[temp_w*4 +:temp_w] = v1115obus[temp_w*1 +:temp_w];
assign v1115ibus[data_w*1 +:data_w] = c251obus[data_w*4 +:data_w];
assign c251ibus[temp_w*5 +:temp_w] = v1403obus[temp_w*1 +:temp_w];
assign v1403ibus[data_w*1 +:data_w] = c251obus[data_w*5 +:data_w];
assign c251ibus[temp_w*6 +:temp_w] = v1499obus[temp_w*0 +:temp_w];
assign v1499ibus[data_w*0 +:data_w] = c251obus[data_w*6 +:data_w];
assign c252ibus[temp_w*0 +:temp_w] = v372obus[temp_w*0 +:temp_w];
assign v372ibus[data_w*0 +:data_w] = c252obus[data_w*0 +:data_w];
assign c252ibus[temp_w*1 +:temp_w] = v466obus[temp_w*0 +:temp_w];
assign v466ibus[data_w*0 +:data_w] = c252obus[data_w*1 +:data_w];
assign c252ibus[temp_w*2 +:temp_w] = v525obus[temp_w*1 +:temp_w];
assign v525ibus[data_w*1 +:data_w] = c252obus[data_w*2 +:data_w];
assign c252ibus[temp_w*3 +:temp_w] = v765obus[temp_w*1 +:temp_w];
assign v765ibus[data_w*1 +:data_w] = c252obus[data_w*3 +:data_w];
assign c252ibus[temp_w*4 +:temp_w] = v1116obus[temp_w*1 +:temp_w];
assign v1116ibus[data_w*1 +:data_w] = c252obus[data_w*4 +:data_w];
assign c252ibus[temp_w*5 +:temp_w] = v1404obus[temp_w*1 +:temp_w];
assign v1404ibus[data_w*1 +:data_w] = c252obus[data_w*5 +:data_w];
assign c252ibus[temp_w*6 +:temp_w] = v1500obus[temp_w*0 +:temp_w];
assign v1500ibus[data_w*0 +:data_w] = c252obus[data_w*6 +:data_w];
assign c253ibus[temp_w*0 +:temp_w] = v373obus[temp_w*0 +:temp_w];
assign v373ibus[data_w*0 +:data_w] = c253obus[data_w*0 +:data_w];
assign c253ibus[temp_w*1 +:temp_w] = v467obus[temp_w*0 +:temp_w];
assign v467ibus[data_w*0 +:data_w] = c253obus[data_w*1 +:data_w];
assign c253ibus[temp_w*2 +:temp_w] = v526obus[temp_w*1 +:temp_w];
assign v526ibus[data_w*1 +:data_w] = c253obus[data_w*2 +:data_w];
assign c253ibus[temp_w*3 +:temp_w] = v766obus[temp_w*1 +:temp_w];
assign v766ibus[data_w*1 +:data_w] = c253obus[data_w*3 +:data_w];
assign c253ibus[temp_w*4 +:temp_w] = v1117obus[temp_w*1 +:temp_w];
assign v1117ibus[data_w*1 +:data_w] = c253obus[data_w*4 +:data_w];
assign c253ibus[temp_w*5 +:temp_w] = v1405obus[temp_w*1 +:temp_w];
assign v1405ibus[data_w*1 +:data_w] = c253obus[data_w*5 +:data_w];
assign c253ibus[temp_w*6 +:temp_w] = v1501obus[temp_w*0 +:temp_w];
assign v1501ibus[data_w*0 +:data_w] = c253obus[data_w*6 +:data_w];
assign c254ibus[temp_w*0 +:temp_w] = v374obus[temp_w*0 +:temp_w];
assign v374ibus[data_w*0 +:data_w] = c254obus[data_w*0 +:data_w];
assign c254ibus[temp_w*1 +:temp_w] = v468obus[temp_w*0 +:temp_w];
assign v468ibus[data_w*0 +:data_w] = c254obus[data_w*1 +:data_w];
assign c254ibus[temp_w*2 +:temp_w] = v527obus[temp_w*1 +:temp_w];
assign v527ibus[data_w*1 +:data_w] = c254obus[data_w*2 +:data_w];
assign c254ibus[temp_w*3 +:temp_w] = v767obus[temp_w*1 +:temp_w];
assign v767ibus[data_w*1 +:data_w] = c254obus[data_w*3 +:data_w];
assign c254ibus[temp_w*4 +:temp_w] = v1118obus[temp_w*1 +:temp_w];
assign v1118ibus[data_w*1 +:data_w] = c254obus[data_w*4 +:data_w];
assign c254ibus[temp_w*5 +:temp_w] = v1406obus[temp_w*1 +:temp_w];
assign v1406ibus[data_w*1 +:data_w] = c254obus[data_w*5 +:data_w];
assign c254ibus[temp_w*6 +:temp_w] = v1502obus[temp_w*0 +:temp_w];
assign v1502ibus[data_w*0 +:data_w] = c254obus[data_w*6 +:data_w];
assign c255ibus[temp_w*0 +:temp_w] = v375obus[temp_w*0 +:temp_w];
assign v375ibus[data_w*0 +:data_w] = c255obus[data_w*0 +:data_w];
assign c255ibus[temp_w*1 +:temp_w] = v469obus[temp_w*0 +:temp_w];
assign v469ibus[data_w*0 +:data_w] = c255obus[data_w*1 +:data_w];
assign c255ibus[temp_w*2 +:temp_w] = v528obus[temp_w*1 +:temp_w];
assign v528ibus[data_w*1 +:data_w] = c255obus[data_w*2 +:data_w];
assign c255ibus[temp_w*3 +:temp_w] = v672obus[temp_w*1 +:temp_w];
assign v672ibus[data_w*1 +:data_w] = c255obus[data_w*3 +:data_w];
assign c255ibus[temp_w*4 +:temp_w] = v1119obus[temp_w*1 +:temp_w];
assign v1119ibus[data_w*1 +:data_w] = c255obus[data_w*4 +:data_w];
assign c255ibus[temp_w*5 +:temp_w] = v1407obus[temp_w*1 +:temp_w];
assign v1407ibus[data_w*1 +:data_w] = c255obus[data_w*5 +:data_w];
assign c255ibus[temp_w*6 +:temp_w] = v1503obus[temp_w*0 +:temp_w];
assign v1503ibus[data_w*0 +:data_w] = c255obus[data_w*6 +:data_w];
assign c256ibus[temp_w*0 +:temp_w] = v376obus[temp_w*0 +:temp_w];
assign v376ibus[data_w*0 +:data_w] = c256obus[data_w*0 +:data_w];
assign c256ibus[temp_w*1 +:temp_w] = v470obus[temp_w*0 +:temp_w];
assign v470ibus[data_w*0 +:data_w] = c256obus[data_w*1 +:data_w];
assign c256ibus[temp_w*2 +:temp_w] = v529obus[temp_w*1 +:temp_w];
assign v529ibus[data_w*1 +:data_w] = c256obus[data_w*2 +:data_w];
assign c256ibus[temp_w*3 +:temp_w] = v673obus[temp_w*1 +:temp_w];
assign v673ibus[data_w*1 +:data_w] = c256obus[data_w*3 +:data_w];
assign c256ibus[temp_w*4 +:temp_w] = v1120obus[temp_w*1 +:temp_w];
assign v1120ibus[data_w*1 +:data_w] = c256obus[data_w*4 +:data_w];
assign c256ibus[temp_w*5 +:temp_w] = v1408obus[temp_w*1 +:temp_w];
assign v1408ibus[data_w*1 +:data_w] = c256obus[data_w*5 +:data_w];
assign c256ibus[temp_w*6 +:temp_w] = v1504obus[temp_w*0 +:temp_w];
assign v1504ibus[data_w*0 +:data_w] = c256obus[data_w*6 +:data_w];
assign c257ibus[temp_w*0 +:temp_w] = v377obus[temp_w*0 +:temp_w];
assign v377ibus[data_w*0 +:data_w] = c257obus[data_w*0 +:data_w];
assign c257ibus[temp_w*1 +:temp_w] = v471obus[temp_w*0 +:temp_w];
assign v471ibus[data_w*0 +:data_w] = c257obus[data_w*1 +:data_w];
assign c257ibus[temp_w*2 +:temp_w] = v530obus[temp_w*1 +:temp_w];
assign v530ibus[data_w*1 +:data_w] = c257obus[data_w*2 +:data_w];
assign c257ibus[temp_w*3 +:temp_w] = v674obus[temp_w*1 +:temp_w];
assign v674ibus[data_w*1 +:data_w] = c257obus[data_w*3 +:data_w];
assign c257ibus[temp_w*4 +:temp_w] = v1121obus[temp_w*1 +:temp_w];
assign v1121ibus[data_w*1 +:data_w] = c257obus[data_w*4 +:data_w];
assign c257ibus[temp_w*5 +:temp_w] = v1409obus[temp_w*1 +:temp_w];
assign v1409ibus[data_w*1 +:data_w] = c257obus[data_w*5 +:data_w];
assign c257ibus[temp_w*6 +:temp_w] = v1505obus[temp_w*0 +:temp_w];
assign v1505ibus[data_w*0 +:data_w] = c257obus[data_w*6 +:data_w];
assign c258ibus[temp_w*0 +:temp_w] = v378obus[temp_w*0 +:temp_w];
assign v378ibus[data_w*0 +:data_w] = c258obus[data_w*0 +:data_w];
assign c258ibus[temp_w*1 +:temp_w] = v472obus[temp_w*0 +:temp_w];
assign v472ibus[data_w*0 +:data_w] = c258obus[data_w*1 +:data_w];
assign c258ibus[temp_w*2 +:temp_w] = v531obus[temp_w*1 +:temp_w];
assign v531ibus[data_w*1 +:data_w] = c258obus[data_w*2 +:data_w];
assign c258ibus[temp_w*3 +:temp_w] = v675obus[temp_w*1 +:temp_w];
assign v675ibus[data_w*1 +:data_w] = c258obus[data_w*3 +:data_w];
assign c258ibus[temp_w*4 +:temp_w] = v1122obus[temp_w*1 +:temp_w];
assign v1122ibus[data_w*1 +:data_w] = c258obus[data_w*4 +:data_w];
assign c258ibus[temp_w*5 +:temp_w] = v1410obus[temp_w*1 +:temp_w];
assign v1410ibus[data_w*1 +:data_w] = c258obus[data_w*5 +:data_w];
assign c258ibus[temp_w*6 +:temp_w] = v1506obus[temp_w*0 +:temp_w];
assign v1506ibus[data_w*0 +:data_w] = c258obus[data_w*6 +:data_w];
assign c259ibus[temp_w*0 +:temp_w] = v379obus[temp_w*0 +:temp_w];
assign v379ibus[data_w*0 +:data_w] = c259obus[data_w*0 +:data_w];
assign c259ibus[temp_w*1 +:temp_w] = v473obus[temp_w*0 +:temp_w];
assign v473ibus[data_w*0 +:data_w] = c259obus[data_w*1 +:data_w];
assign c259ibus[temp_w*2 +:temp_w] = v532obus[temp_w*1 +:temp_w];
assign v532ibus[data_w*1 +:data_w] = c259obus[data_w*2 +:data_w];
assign c259ibus[temp_w*3 +:temp_w] = v676obus[temp_w*1 +:temp_w];
assign v676ibus[data_w*1 +:data_w] = c259obus[data_w*3 +:data_w];
assign c259ibus[temp_w*4 +:temp_w] = v1123obus[temp_w*1 +:temp_w];
assign v1123ibus[data_w*1 +:data_w] = c259obus[data_w*4 +:data_w];
assign c259ibus[temp_w*5 +:temp_w] = v1411obus[temp_w*1 +:temp_w];
assign v1411ibus[data_w*1 +:data_w] = c259obus[data_w*5 +:data_w];
assign c259ibus[temp_w*6 +:temp_w] = v1507obus[temp_w*0 +:temp_w];
assign v1507ibus[data_w*0 +:data_w] = c259obus[data_w*6 +:data_w];
assign c260ibus[temp_w*0 +:temp_w] = v380obus[temp_w*0 +:temp_w];
assign v380ibus[data_w*0 +:data_w] = c260obus[data_w*0 +:data_w];
assign c260ibus[temp_w*1 +:temp_w] = v474obus[temp_w*0 +:temp_w];
assign v474ibus[data_w*0 +:data_w] = c260obus[data_w*1 +:data_w];
assign c260ibus[temp_w*2 +:temp_w] = v533obus[temp_w*1 +:temp_w];
assign v533ibus[data_w*1 +:data_w] = c260obus[data_w*2 +:data_w];
assign c260ibus[temp_w*3 +:temp_w] = v677obus[temp_w*1 +:temp_w];
assign v677ibus[data_w*1 +:data_w] = c260obus[data_w*3 +:data_w];
assign c260ibus[temp_w*4 +:temp_w] = v1124obus[temp_w*1 +:temp_w];
assign v1124ibus[data_w*1 +:data_w] = c260obus[data_w*4 +:data_w];
assign c260ibus[temp_w*5 +:temp_w] = v1412obus[temp_w*1 +:temp_w];
assign v1412ibus[data_w*1 +:data_w] = c260obus[data_w*5 +:data_w];
assign c260ibus[temp_w*6 +:temp_w] = v1508obus[temp_w*0 +:temp_w];
assign v1508ibus[data_w*0 +:data_w] = c260obus[data_w*6 +:data_w];
assign c261ibus[temp_w*0 +:temp_w] = v381obus[temp_w*0 +:temp_w];
assign v381ibus[data_w*0 +:data_w] = c261obus[data_w*0 +:data_w];
assign c261ibus[temp_w*1 +:temp_w] = v475obus[temp_w*0 +:temp_w];
assign v475ibus[data_w*0 +:data_w] = c261obus[data_w*1 +:data_w];
assign c261ibus[temp_w*2 +:temp_w] = v534obus[temp_w*1 +:temp_w];
assign v534ibus[data_w*1 +:data_w] = c261obus[data_w*2 +:data_w];
assign c261ibus[temp_w*3 +:temp_w] = v678obus[temp_w*1 +:temp_w];
assign v678ibus[data_w*1 +:data_w] = c261obus[data_w*3 +:data_w];
assign c261ibus[temp_w*4 +:temp_w] = v1125obus[temp_w*1 +:temp_w];
assign v1125ibus[data_w*1 +:data_w] = c261obus[data_w*4 +:data_w];
assign c261ibus[temp_w*5 +:temp_w] = v1413obus[temp_w*1 +:temp_w];
assign v1413ibus[data_w*1 +:data_w] = c261obus[data_w*5 +:data_w];
assign c261ibus[temp_w*6 +:temp_w] = v1509obus[temp_w*0 +:temp_w];
assign v1509ibus[data_w*0 +:data_w] = c261obus[data_w*6 +:data_w];
assign c262ibus[temp_w*0 +:temp_w] = v382obus[temp_w*0 +:temp_w];
assign v382ibus[data_w*0 +:data_w] = c262obus[data_w*0 +:data_w];
assign c262ibus[temp_w*1 +:temp_w] = v476obus[temp_w*0 +:temp_w];
assign v476ibus[data_w*0 +:data_w] = c262obus[data_w*1 +:data_w];
assign c262ibus[temp_w*2 +:temp_w] = v535obus[temp_w*1 +:temp_w];
assign v535ibus[data_w*1 +:data_w] = c262obus[data_w*2 +:data_w];
assign c262ibus[temp_w*3 +:temp_w] = v679obus[temp_w*1 +:temp_w];
assign v679ibus[data_w*1 +:data_w] = c262obus[data_w*3 +:data_w];
assign c262ibus[temp_w*4 +:temp_w] = v1126obus[temp_w*1 +:temp_w];
assign v1126ibus[data_w*1 +:data_w] = c262obus[data_w*4 +:data_w];
assign c262ibus[temp_w*5 +:temp_w] = v1414obus[temp_w*1 +:temp_w];
assign v1414ibus[data_w*1 +:data_w] = c262obus[data_w*5 +:data_w];
assign c262ibus[temp_w*6 +:temp_w] = v1510obus[temp_w*0 +:temp_w];
assign v1510ibus[data_w*0 +:data_w] = c262obus[data_w*6 +:data_w];
assign c263ibus[temp_w*0 +:temp_w] = v383obus[temp_w*0 +:temp_w];
assign v383ibus[data_w*0 +:data_w] = c263obus[data_w*0 +:data_w];
assign c263ibus[temp_w*1 +:temp_w] = v477obus[temp_w*0 +:temp_w];
assign v477ibus[data_w*0 +:data_w] = c263obus[data_w*1 +:data_w];
assign c263ibus[temp_w*2 +:temp_w] = v536obus[temp_w*1 +:temp_w];
assign v536ibus[data_w*1 +:data_w] = c263obus[data_w*2 +:data_w];
assign c263ibus[temp_w*3 +:temp_w] = v680obus[temp_w*1 +:temp_w];
assign v680ibus[data_w*1 +:data_w] = c263obus[data_w*3 +:data_w];
assign c263ibus[temp_w*4 +:temp_w] = v1127obus[temp_w*1 +:temp_w];
assign v1127ibus[data_w*1 +:data_w] = c263obus[data_w*4 +:data_w];
assign c263ibus[temp_w*5 +:temp_w] = v1415obus[temp_w*1 +:temp_w];
assign v1415ibus[data_w*1 +:data_w] = c263obus[data_w*5 +:data_w];
assign c263ibus[temp_w*6 +:temp_w] = v1511obus[temp_w*0 +:temp_w];
assign v1511ibus[data_w*0 +:data_w] = c263obus[data_w*6 +:data_w];
assign c264ibus[temp_w*0 +:temp_w] = v288obus[temp_w*0 +:temp_w];
assign v288ibus[data_w*0 +:data_w] = c264obus[data_w*0 +:data_w];
assign c264ibus[temp_w*1 +:temp_w] = v478obus[temp_w*0 +:temp_w];
assign v478ibus[data_w*0 +:data_w] = c264obus[data_w*1 +:data_w];
assign c264ibus[temp_w*2 +:temp_w] = v537obus[temp_w*1 +:temp_w];
assign v537ibus[data_w*1 +:data_w] = c264obus[data_w*2 +:data_w];
assign c264ibus[temp_w*3 +:temp_w] = v681obus[temp_w*1 +:temp_w];
assign v681ibus[data_w*1 +:data_w] = c264obus[data_w*3 +:data_w];
assign c264ibus[temp_w*4 +:temp_w] = v1128obus[temp_w*1 +:temp_w];
assign v1128ibus[data_w*1 +:data_w] = c264obus[data_w*4 +:data_w];
assign c264ibus[temp_w*5 +:temp_w] = v1416obus[temp_w*1 +:temp_w];
assign v1416ibus[data_w*1 +:data_w] = c264obus[data_w*5 +:data_w];
assign c264ibus[temp_w*6 +:temp_w] = v1512obus[temp_w*0 +:temp_w];
assign v1512ibus[data_w*0 +:data_w] = c264obus[data_w*6 +:data_w];
assign c265ibus[temp_w*0 +:temp_w] = v289obus[temp_w*0 +:temp_w];
assign v289ibus[data_w*0 +:data_w] = c265obus[data_w*0 +:data_w];
assign c265ibus[temp_w*1 +:temp_w] = v479obus[temp_w*0 +:temp_w];
assign v479ibus[data_w*0 +:data_w] = c265obus[data_w*1 +:data_w];
assign c265ibus[temp_w*2 +:temp_w] = v538obus[temp_w*1 +:temp_w];
assign v538ibus[data_w*1 +:data_w] = c265obus[data_w*2 +:data_w];
assign c265ibus[temp_w*3 +:temp_w] = v682obus[temp_w*1 +:temp_w];
assign v682ibus[data_w*1 +:data_w] = c265obus[data_w*3 +:data_w];
assign c265ibus[temp_w*4 +:temp_w] = v1129obus[temp_w*1 +:temp_w];
assign v1129ibus[data_w*1 +:data_w] = c265obus[data_w*4 +:data_w];
assign c265ibus[temp_w*5 +:temp_w] = v1417obus[temp_w*1 +:temp_w];
assign v1417ibus[data_w*1 +:data_w] = c265obus[data_w*5 +:data_w];
assign c265ibus[temp_w*6 +:temp_w] = v1513obus[temp_w*0 +:temp_w];
assign v1513ibus[data_w*0 +:data_w] = c265obus[data_w*6 +:data_w];
assign c266ibus[temp_w*0 +:temp_w] = v290obus[temp_w*0 +:temp_w];
assign v290ibus[data_w*0 +:data_w] = c266obus[data_w*0 +:data_w];
assign c266ibus[temp_w*1 +:temp_w] = v384obus[temp_w*0 +:temp_w];
assign v384ibus[data_w*0 +:data_w] = c266obus[data_w*1 +:data_w];
assign c266ibus[temp_w*2 +:temp_w] = v539obus[temp_w*1 +:temp_w];
assign v539ibus[data_w*1 +:data_w] = c266obus[data_w*2 +:data_w];
assign c266ibus[temp_w*3 +:temp_w] = v683obus[temp_w*1 +:temp_w];
assign v683ibus[data_w*1 +:data_w] = c266obus[data_w*3 +:data_w];
assign c266ibus[temp_w*4 +:temp_w] = v1130obus[temp_w*1 +:temp_w];
assign v1130ibus[data_w*1 +:data_w] = c266obus[data_w*4 +:data_w];
assign c266ibus[temp_w*5 +:temp_w] = v1418obus[temp_w*1 +:temp_w];
assign v1418ibus[data_w*1 +:data_w] = c266obus[data_w*5 +:data_w];
assign c266ibus[temp_w*6 +:temp_w] = v1514obus[temp_w*0 +:temp_w];
assign v1514ibus[data_w*0 +:data_w] = c266obus[data_w*6 +:data_w];
assign c267ibus[temp_w*0 +:temp_w] = v291obus[temp_w*0 +:temp_w];
assign v291ibus[data_w*0 +:data_w] = c267obus[data_w*0 +:data_w];
assign c267ibus[temp_w*1 +:temp_w] = v385obus[temp_w*0 +:temp_w];
assign v385ibus[data_w*0 +:data_w] = c267obus[data_w*1 +:data_w];
assign c267ibus[temp_w*2 +:temp_w] = v540obus[temp_w*1 +:temp_w];
assign v540ibus[data_w*1 +:data_w] = c267obus[data_w*2 +:data_w];
assign c267ibus[temp_w*3 +:temp_w] = v684obus[temp_w*1 +:temp_w];
assign v684ibus[data_w*1 +:data_w] = c267obus[data_w*3 +:data_w];
assign c267ibus[temp_w*4 +:temp_w] = v1131obus[temp_w*1 +:temp_w];
assign v1131ibus[data_w*1 +:data_w] = c267obus[data_w*4 +:data_w];
assign c267ibus[temp_w*5 +:temp_w] = v1419obus[temp_w*1 +:temp_w];
assign v1419ibus[data_w*1 +:data_w] = c267obus[data_w*5 +:data_w];
assign c267ibus[temp_w*6 +:temp_w] = v1515obus[temp_w*0 +:temp_w];
assign v1515ibus[data_w*0 +:data_w] = c267obus[data_w*6 +:data_w];
assign c268ibus[temp_w*0 +:temp_w] = v292obus[temp_w*0 +:temp_w];
assign v292ibus[data_w*0 +:data_w] = c268obus[data_w*0 +:data_w];
assign c268ibus[temp_w*1 +:temp_w] = v386obus[temp_w*0 +:temp_w];
assign v386ibus[data_w*0 +:data_w] = c268obus[data_w*1 +:data_w];
assign c268ibus[temp_w*2 +:temp_w] = v541obus[temp_w*1 +:temp_w];
assign v541ibus[data_w*1 +:data_w] = c268obus[data_w*2 +:data_w];
assign c268ibus[temp_w*3 +:temp_w] = v685obus[temp_w*1 +:temp_w];
assign v685ibus[data_w*1 +:data_w] = c268obus[data_w*3 +:data_w];
assign c268ibus[temp_w*4 +:temp_w] = v1132obus[temp_w*1 +:temp_w];
assign v1132ibus[data_w*1 +:data_w] = c268obus[data_w*4 +:data_w];
assign c268ibus[temp_w*5 +:temp_w] = v1420obus[temp_w*1 +:temp_w];
assign v1420ibus[data_w*1 +:data_w] = c268obus[data_w*5 +:data_w];
assign c268ibus[temp_w*6 +:temp_w] = v1516obus[temp_w*0 +:temp_w];
assign v1516ibus[data_w*0 +:data_w] = c268obus[data_w*6 +:data_w];
assign c269ibus[temp_w*0 +:temp_w] = v293obus[temp_w*0 +:temp_w];
assign v293ibus[data_w*0 +:data_w] = c269obus[data_w*0 +:data_w];
assign c269ibus[temp_w*1 +:temp_w] = v387obus[temp_w*0 +:temp_w];
assign v387ibus[data_w*0 +:data_w] = c269obus[data_w*1 +:data_w];
assign c269ibus[temp_w*2 +:temp_w] = v542obus[temp_w*1 +:temp_w];
assign v542ibus[data_w*1 +:data_w] = c269obus[data_w*2 +:data_w];
assign c269ibus[temp_w*3 +:temp_w] = v686obus[temp_w*1 +:temp_w];
assign v686ibus[data_w*1 +:data_w] = c269obus[data_w*3 +:data_w];
assign c269ibus[temp_w*4 +:temp_w] = v1133obus[temp_w*1 +:temp_w];
assign v1133ibus[data_w*1 +:data_w] = c269obus[data_w*4 +:data_w];
assign c269ibus[temp_w*5 +:temp_w] = v1421obus[temp_w*1 +:temp_w];
assign v1421ibus[data_w*1 +:data_w] = c269obus[data_w*5 +:data_w];
assign c269ibus[temp_w*6 +:temp_w] = v1517obus[temp_w*0 +:temp_w];
assign v1517ibus[data_w*0 +:data_w] = c269obus[data_w*6 +:data_w];
assign c270ibus[temp_w*0 +:temp_w] = v294obus[temp_w*0 +:temp_w];
assign v294ibus[data_w*0 +:data_w] = c270obus[data_w*0 +:data_w];
assign c270ibus[temp_w*1 +:temp_w] = v388obus[temp_w*0 +:temp_w];
assign v388ibus[data_w*0 +:data_w] = c270obus[data_w*1 +:data_w];
assign c270ibus[temp_w*2 +:temp_w] = v543obus[temp_w*1 +:temp_w];
assign v543ibus[data_w*1 +:data_w] = c270obus[data_w*2 +:data_w];
assign c270ibus[temp_w*3 +:temp_w] = v687obus[temp_w*1 +:temp_w];
assign v687ibus[data_w*1 +:data_w] = c270obus[data_w*3 +:data_w];
assign c270ibus[temp_w*4 +:temp_w] = v1134obus[temp_w*1 +:temp_w];
assign v1134ibus[data_w*1 +:data_w] = c270obus[data_w*4 +:data_w];
assign c270ibus[temp_w*5 +:temp_w] = v1422obus[temp_w*1 +:temp_w];
assign v1422ibus[data_w*1 +:data_w] = c270obus[data_w*5 +:data_w];
assign c270ibus[temp_w*6 +:temp_w] = v1518obus[temp_w*0 +:temp_w];
assign v1518ibus[data_w*0 +:data_w] = c270obus[data_w*6 +:data_w];
assign c271ibus[temp_w*0 +:temp_w] = v295obus[temp_w*0 +:temp_w];
assign v295ibus[data_w*0 +:data_w] = c271obus[data_w*0 +:data_w];
assign c271ibus[temp_w*1 +:temp_w] = v389obus[temp_w*0 +:temp_w];
assign v389ibus[data_w*0 +:data_w] = c271obus[data_w*1 +:data_w];
assign c271ibus[temp_w*2 +:temp_w] = v544obus[temp_w*1 +:temp_w];
assign v544ibus[data_w*1 +:data_w] = c271obus[data_w*2 +:data_w];
assign c271ibus[temp_w*3 +:temp_w] = v688obus[temp_w*1 +:temp_w];
assign v688ibus[data_w*1 +:data_w] = c271obus[data_w*3 +:data_w];
assign c271ibus[temp_w*4 +:temp_w] = v1135obus[temp_w*1 +:temp_w];
assign v1135ibus[data_w*1 +:data_w] = c271obus[data_w*4 +:data_w];
assign c271ibus[temp_w*5 +:temp_w] = v1423obus[temp_w*1 +:temp_w];
assign v1423ibus[data_w*1 +:data_w] = c271obus[data_w*5 +:data_w];
assign c271ibus[temp_w*6 +:temp_w] = v1519obus[temp_w*0 +:temp_w];
assign v1519ibus[data_w*0 +:data_w] = c271obus[data_w*6 +:data_w];
assign c272ibus[temp_w*0 +:temp_w] = v296obus[temp_w*0 +:temp_w];
assign v296ibus[data_w*0 +:data_w] = c272obus[data_w*0 +:data_w];
assign c272ibus[temp_w*1 +:temp_w] = v390obus[temp_w*0 +:temp_w];
assign v390ibus[data_w*0 +:data_w] = c272obus[data_w*1 +:data_w];
assign c272ibus[temp_w*2 +:temp_w] = v545obus[temp_w*1 +:temp_w];
assign v545ibus[data_w*1 +:data_w] = c272obus[data_w*2 +:data_w];
assign c272ibus[temp_w*3 +:temp_w] = v689obus[temp_w*1 +:temp_w];
assign v689ibus[data_w*1 +:data_w] = c272obus[data_w*3 +:data_w];
assign c272ibus[temp_w*4 +:temp_w] = v1136obus[temp_w*1 +:temp_w];
assign v1136ibus[data_w*1 +:data_w] = c272obus[data_w*4 +:data_w];
assign c272ibus[temp_w*5 +:temp_w] = v1424obus[temp_w*1 +:temp_w];
assign v1424ibus[data_w*1 +:data_w] = c272obus[data_w*5 +:data_w];
assign c272ibus[temp_w*6 +:temp_w] = v1520obus[temp_w*0 +:temp_w];
assign v1520ibus[data_w*0 +:data_w] = c272obus[data_w*6 +:data_w];
assign c273ibus[temp_w*0 +:temp_w] = v297obus[temp_w*0 +:temp_w];
assign v297ibus[data_w*0 +:data_w] = c273obus[data_w*0 +:data_w];
assign c273ibus[temp_w*1 +:temp_w] = v391obus[temp_w*0 +:temp_w];
assign v391ibus[data_w*0 +:data_w] = c273obus[data_w*1 +:data_w];
assign c273ibus[temp_w*2 +:temp_w] = v546obus[temp_w*1 +:temp_w];
assign v546ibus[data_w*1 +:data_w] = c273obus[data_w*2 +:data_w];
assign c273ibus[temp_w*3 +:temp_w] = v690obus[temp_w*1 +:temp_w];
assign v690ibus[data_w*1 +:data_w] = c273obus[data_w*3 +:data_w];
assign c273ibus[temp_w*4 +:temp_w] = v1137obus[temp_w*1 +:temp_w];
assign v1137ibus[data_w*1 +:data_w] = c273obus[data_w*4 +:data_w];
assign c273ibus[temp_w*5 +:temp_w] = v1425obus[temp_w*1 +:temp_w];
assign v1425ibus[data_w*1 +:data_w] = c273obus[data_w*5 +:data_w];
assign c273ibus[temp_w*6 +:temp_w] = v1521obus[temp_w*0 +:temp_w];
assign v1521ibus[data_w*0 +:data_w] = c273obus[data_w*6 +:data_w];
assign c274ibus[temp_w*0 +:temp_w] = v298obus[temp_w*0 +:temp_w];
assign v298ibus[data_w*0 +:data_w] = c274obus[data_w*0 +:data_w];
assign c274ibus[temp_w*1 +:temp_w] = v392obus[temp_w*0 +:temp_w];
assign v392ibus[data_w*0 +:data_w] = c274obus[data_w*1 +:data_w];
assign c274ibus[temp_w*2 +:temp_w] = v547obus[temp_w*1 +:temp_w];
assign v547ibus[data_w*1 +:data_w] = c274obus[data_w*2 +:data_w];
assign c274ibus[temp_w*3 +:temp_w] = v691obus[temp_w*1 +:temp_w];
assign v691ibus[data_w*1 +:data_w] = c274obus[data_w*3 +:data_w];
assign c274ibus[temp_w*4 +:temp_w] = v1138obus[temp_w*1 +:temp_w];
assign v1138ibus[data_w*1 +:data_w] = c274obus[data_w*4 +:data_w];
assign c274ibus[temp_w*5 +:temp_w] = v1426obus[temp_w*1 +:temp_w];
assign v1426ibus[data_w*1 +:data_w] = c274obus[data_w*5 +:data_w];
assign c274ibus[temp_w*6 +:temp_w] = v1522obus[temp_w*0 +:temp_w];
assign v1522ibus[data_w*0 +:data_w] = c274obus[data_w*6 +:data_w];
assign c275ibus[temp_w*0 +:temp_w] = v299obus[temp_w*0 +:temp_w];
assign v299ibus[data_w*0 +:data_w] = c275obus[data_w*0 +:data_w];
assign c275ibus[temp_w*1 +:temp_w] = v393obus[temp_w*0 +:temp_w];
assign v393ibus[data_w*0 +:data_w] = c275obus[data_w*1 +:data_w];
assign c275ibus[temp_w*2 +:temp_w] = v548obus[temp_w*1 +:temp_w];
assign v548ibus[data_w*1 +:data_w] = c275obus[data_w*2 +:data_w];
assign c275ibus[temp_w*3 +:temp_w] = v692obus[temp_w*1 +:temp_w];
assign v692ibus[data_w*1 +:data_w] = c275obus[data_w*3 +:data_w];
assign c275ibus[temp_w*4 +:temp_w] = v1139obus[temp_w*1 +:temp_w];
assign v1139ibus[data_w*1 +:data_w] = c275obus[data_w*4 +:data_w];
assign c275ibus[temp_w*5 +:temp_w] = v1427obus[temp_w*1 +:temp_w];
assign v1427ibus[data_w*1 +:data_w] = c275obus[data_w*5 +:data_w];
assign c275ibus[temp_w*6 +:temp_w] = v1523obus[temp_w*0 +:temp_w];
assign v1523ibus[data_w*0 +:data_w] = c275obus[data_w*6 +:data_w];
assign c276ibus[temp_w*0 +:temp_w] = v300obus[temp_w*0 +:temp_w];
assign v300ibus[data_w*0 +:data_w] = c276obus[data_w*0 +:data_w];
assign c276ibus[temp_w*1 +:temp_w] = v394obus[temp_w*0 +:temp_w];
assign v394ibus[data_w*0 +:data_w] = c276obus[data_w*1 +:data_w];
assign c276ibus[temp_w*2 +:temp_w] = v549obus[temp_w*1 +:temp_w];
assign v549ibus[data_w*1 +:data_w] = c276obus[data_w*2 +:data_w];
assign c276ibus[temp_w*3 +:temp_w] = v693obus[temp_w*1 +:temp_w];
assign v693ibus[data_w*1 +:data_w] = c276obus[data_w*3 +:data_w];
assign c276ibus[temp_w*4 +:temp_w] = v1140obus[temp_w*1 +:temp_w];
assign v1140ibus[data_w*1 +:data_w] = c276obus[data_w*4 +:data_w];
assign c276ibus[temp_w*5 +:temp_w] = v1428obus[temp_w*1 +:temp_w];
assign v1428ibus[data_w*1 +:data_w] = c276obus[data_w*5 +:data_w];
assign c276ibus[temp_w*6 +:temp_w] = v1524obus[temp_w*0 +:temp_w];
assign v1524ibus[data_w*0 +:data_w] = c276obus[data_w*6 +:data_w];
assign c277ibus[temp_w*0 +:temp_w] = v301obus[temp_w*0 +:temp_w];
assign v301ibus[data_w*0 +:data_w] = c277obus[data_w*0 +:data_w];
assign c277ibus[temp_w*1 +:temp_w] = v395obus[temp_w*0 +:temp_w];
assign v395ibus[data_w*0 +:data_w] = c277obus[data_w*1 +:data_w];
assign c277ibus[temp_w*2 +:temp_w] = v550obus[temp_w*1 +:temp_w];
assign v550ibus[data_w*1 +:data_w] = c277obus[data_w*2 +:data_w];
assign c277ibus[temp_w*3 +:temp_w] = v694obus[temp_w*1 +:temp_w];
assign v694ibus[data_w*1 +:data_w] = c277obus[data_w*3 +:data_w];
assign c277ibus[temp_w*4 +:temp_w] = v1141obus[temp_w*1 +:temp_w];
assign v1141ibus[data_w*1 +:data_w] = c277obus[data_w*4 +:data_w];
assign c277ibus[temp_w*5 +:temp_w] = v1429obus[temp_w*1 +:temp_w];
assign v1429ibus[data_w*1 +:data_w] = c277obus[data_w*5 +:data_w];
assign c277ibus[temp_w*6 +:temp_w] = v1525obus[temp_w*0 +:temp_w];
assign v1525ibus[data_w*0 +:data_w] = c277obus[data_w*6 +:data_w];
assign c278ibus[temp_w*0 +:temp_w] = v302obus[temp_w*0 +:temp_w];
assign v302ibus[data_w*0 +:data_w] = c278obus[data_w*0 +:data_w];
assign c278ibus[temp_w*1 +:temp_w] = v396obus[temp_w*0 +:temp_w];
assign v396ibus[data_w*0 +:data_w] = c278obus[data_w*1 +:data_w];
assign c278ibus[temp_w*2 +:temp_w] = v551obus[temp_w*1 +:temp_w];
assign v551ibus[data_w*1 +:data_w] = c278obus[data_w*2 +:data_w];
assign c278ibus[temp_w*3 +:temp_w] = v695obus[temp_w*1 +:temp_w];
assign v695ibus[data_w*1 +:data_w] = c278obus[data_w*3 +:data_w];
assign c278ibus[temp_w*4 +:temp_w] = v1142obus[temp_w*1 +:temp_w];
assign v1142ibus[data_w*1 +:data_w] = c278obus[data_w*4 +:data_w];
assign c278ibus[temp_w*5 +:temp_w] = v1430obus[temp_w*1 +:temp_w];
assign v1430ibus[data_w*1 +:data_w] = c278obus[data_w*5 +:data_w];
assign c278ibus[temp_w*6 +:temp_w] = v1526obus[temp_w*0 +:temp_w];
assign v1526ibus[data_w*0 +:data_w] = c278obus[data_w*6 +:data_w];
assign c279ibus[temp_w*0 +:temp_w] = v303obus[temp_w*0 +:temp_w];
assign v303ibus[data_w*0 +:data_w] = c279obus[data_w*0 +:data_w];
assign c279ibus[temp_w*1 +:temp_w] = v397obus[temp_w*0 +:temp_w];
assign v397ibus[data_w*0 +:data_w] = c279obus[data_w*1 +:data_w];
assign c279ibus[temp_w*2 +:temp_w] = v552obus[temp_w*1 +:temp_w];
assign v552ibus[data_w*1 +:data_w] = c279obus[data_w*2 +:data_w];
assign c279ibus[temp_w*3 +:temp_w] = v696obus[temp_w*1 +:temp_w];
assign v696ibus[data_w*1 +:data_w] = c279obus[data_w*3 +:data_w];
assign c279ibus[temp_w*4 +:temp_w] = v1143obus[temp_w*1 +:temp_w];
assign v1143ibus[data_w*1 +:data_w] = c279obus[data_w*4 +:data_w];
assign c279ibus[temp_w*5 +:temp_w] = v1431obus[temp_w*1 +:temp_w];
assign v1431ibus[data_w*1 +:data_w] = c279obus[data_w*5 +:data_w];
assign c279ibus[temp_w*6 +:temp_w] = v1527obus[temp_w*0 +:temp_w];
assign v1527ibus[data_w*0 +:data_w] = c279obus[data_w*6 +:data_w];
assign c280ibus[temp_w*0 +:temp_w] = v304obus[temp_w*0 +:temp_w];
assign v304ibus[data_w*0 +:data_w] = c280obus[data_w*0 +:data_w];
assign c280ibus[temp_w*1 +:temp_w] = v398obus[temp_w*0 +:temp_w];
assign v398ibus[data_w*0 +:data_w] = c280obus[data_w*1 +:data_w];
assign c280ibus[temp_w*2 +:temp_w] = v553obus[temp_w*1 +:temp_w];
assign v553ibus[data_w*1 +:data_w] = c280obus[data_w*2 +:data_w];
assign c280ibus[temp_w*3 +:temp_w] = v697obus[temp_w*1 +:temp_w];
assign v697ibus[data_w*1 +:data_w] = c280obus[data_w*3 +:data_w];
assign c280ibus[temp_w*4 +:temp_w] = v1144obus[temp_w*1 +:temp_w];
assign v1144ibus[data_w*1 +:data_w] = c280obus[data_w*4 +:data_w];
assign c280ibus[temp_w*5 +:temp_w] = v1432obus[temp_w*1 +:temp_w];
assign v1432ibus[data_w*1 +:data_w] = c280obus[data_w*5 +:data_w];
assign c280ibus[temp_w*6 +:temp_w] = v1528obus[temp_w*0 +:temp_w];
assign v1528ibus[data_w*0 +:data_w] = c280obus[data_w*6 +:data_w];
assign c281ibus[temp_w*0 +:temp_w] = v305obus[temp_w*0 +:temp_w];
assign v305ibus[data_w*0 +:data_w] = c281obus[data_w*0 +:data_w];
assign c281ibus[temp_w*1 +:temp_w] = v399obus[temp_w*0 +:temp_w];
assign v399ibus[data_w*0 +:data_w] = c281obus[data_w*1 +:data_w];
assign c281ibus[temp_w*2 +:temp_w] = v554obus[temp_w*1 +:temp_w];
assign v554ibus[data_w*1 +:data_w] = c281obus[data_w*2 +:data_w];
assign c281ibus[temp_w*3 +:temp_w] = v698obus[temp_w*1 +:temp_w];
assign v698ibus[data_w*1 +:data_w] = c281obus[data_w*3 +:data_w];
assign c281ibus[temp_w*4 +:temp_w] = v1145obus[temp_w*1 +:temp_w];
assign v1145ibus[data_w*1 +:data_w] = c281obus[data_w*4 +:data_w];
assign c281ibus[temp_w*5 +:temp_w] = v1433obus[temp_w*1 +:temp_w];
assign v1433ibus[data_w*1 +:data_w] = c281obus[data_w*5 +:data_w];
assign c281ibus[temp_w*6 +:temp_w] = v1529obus[temp_w*0 +:temp_w];
assign v1529ibus[data_w*0 +:data_w] = c281obus[data_w*6 +:data_w];
assign c282ibus[temp_w*0 +:temp_w] = v306obus[temp_w*0 +:temp_w];
assign v306ibus[data_w*0 +:data_w] = c282obus[data_w*0 +:data_w];
assign c282ibus[temp_w*1 +:temp_w] = v400obus[temp_w*0 +:temp_w];
assign v400ibus[data_w*0 +:data_w] = c282obus[data_w*1 +:data_w];
assign c282ibus[temp_w*2 +:temp_w] = v555obus[temp_w*1 +:temp_w];
assign v555ibus[data_w*1 +:data_w] = c282obus[data_w*2 +:data_w];
assign c282ibus[temp_w*3 +:temp_w] = v699obus[temp_w*1 +:temp_w];
assign v699ibus[data_w*1 +:data_w] = c282obus[data_w*3 +:data_w];
assign c282ibus[temp_w*4 +:temp_w] = v1146obus[temp_w*1 +:temp_w];
assign v1146ibus[data_w*1 +:data_w] = c282obus[data_w*4 +:data_w];
assign c282ibus[temp_w*5 +:temp_w] = v1434obus[temp_w*1 +:temp_w];
assign v1434ibus[data_w*1 +:data_w] = c282obus[data_w*5 +:data_w];
assign c282ibus[temp_w*6 +:temp_w] = v1530obus[temp_w*0 +:temp_w];
assign v1530ibus[data_w*0 +:data_w] = c282obus[data_w*6 +:data_w];
assign c283ibus[temp_w*0 +:temp_w] = v307obus[temp_w*0 +:temp_w];
assign v307ibus[data_w*0 +:data_w] = c283obus[data_w*0 +:data_w];
assign c283ibus[temp_w*1 +:temp_w] = v401obus[temp_w*0 +:temp_w];
assign v401ibus[data_w*0 +:data_w] = c283obus[data_w*1 +:data_w];
assign c283ibus[temp_w*2 +:temp_w] = v556obus[temp_w*1 +:temp_w];
assign v556ibus[data_w*1 +:data_w] = c283obus[data_w*2 +:data_w];
assign c283ibus[temp_w*3 +:temp_w] = v700obus[temp_w*1 +:temp_w];
assign v700ibus[data_w*1 +:data_w] = c283obus[data_w*3 +:data_w];
assign c283ibus[temp_w*4 +:temp_w] = v1147obus[temp_w*1 +:temp_w];
assign v1147ibus[data_w*1 +:data_w] = c283obus[data_w*4 +:data_w];
assign c283ibus[temp_w*5 +:temp_w] = v1435obus[temp_w*1 +:temp_w];
assign v1435ibus[data_w*1 +:data_w] = c283obus[data_w*5 +:data_w];
assign c283ibus[temp_w*6 +:temp_w] = v1531obus[temp_w*0 +:temp_w];
assign v1531ibus[data_w*0 +:data_w] = c283obus[data_w*6 +:data_w];
assign c284ibus[temp_w*0 +:temp_w] = v308obus[temp_w*0 +:temp_w];
assign v308ibus[data_w*0 +:data_w] = c284obus[data_w*0 +:data_w];
assign c284ibus[temp_w*1 +:temp_w] = v402obus[temp_w*0 +:temp_w];
assign v402ibus[data_w*0 +:data_w] = c284obus[data_w*1 +:data_w];
assign c284ibus[temp_w*2 +:temp_w] = v557obus[temp_w*1 +:temp_w];
assign v557ibus[data_w*1 +:data_w] = c284obus[data_w*2 +:data_w];
assign c284ibus[temp_w*3 +:temp_w] = v701obus[temp_w*1 +:temp_w];
assign v701ibus[data_w*1 +:data_w] = c284obus[data_w*3 +:data_w];
assign c284ibus[temp_w*4 +:temp_w] = v1148obus[temp_w*1 +:temp_w];
assign v1148ibus[data_w*1 +:data_w] = c284obus[data_w*4 +:data_w];
assign c284ibus[temp_w*5 +:temp_w] = v1436obus[temp_w*1 +:temp_w];
assign v1436ibus[data_w*1 +:data_w] = c284obus[data_w*5 +:data_w];
assign c284ibus[temp_w*6 +:temp_w] = v1532obus[temp_w*0 +:temp_w];
assign v1532ibus[data_w*0 +:data_w] = c284obus[data_w*6 +:data_w];
assign c285ibus[temp_w*0 +:temp_w] = v309obus[temp_w*0 +:temp_w];
assign v309ibus[data_w*0 +:data_w] = c285obus[data_w*0 +:data_w];
assign c285ibus[temp_w*1 +:temp_w] = v403obus[temp_w*0 +:temp_w];
assign v403ibus[data_w*0 +:data_w] = c285obus[data_w*1 +:data_w];
assign c285ibus[temp_w*2 +:temp_w] = v558obus[temp_w*1 +:temp_w];
assign v558ibus[data_w*1 +:data_w] = c285obus[data_w*2 +:data_w];
assign c285ibus[temp_w*3 +:temp_w] = v702obus[temp_w*1 +:temp_w];
assign v702ibus[data_w*1 +:data_w] = c285obus[data_w*3 +:data_w];
assign c285ibus[temp_w*4 +:temp_w] = v1149obus[temp_w*1 +:temp_w];
assign v1149ibus[data_w*1 +:data_w] = c285obus[data_w*4 +:data_w];
assign c285ibus[temp_w*5 +:temp_w] = v1437obus[temp_w*1 +:temp_w];
assign v1437ibus[data_w*1 +:data_w] = c285obus[data_w*5 +:data_w];
assign c285ibus[temp_w*6 +:temp_w] = v1533obus[temp_w*0 +:temp_w];
assign v1533ibus[data_w*0 +:data_w] = c285obus[data_w*6 +:data_w];
assign c286ibus[temp_w*0 +:temp_w] = v310obus[temp_w*0 +:temp_w];
assign v310ibus[data_w*0 +:data_w] = c286obus[data_w*0 +:data_w];
assign c286ibus[temp_w*1 +:temp_w] = v404obus[temp_w*0 +:temp_w];
assign v404ibus[data_w*0 +:data_w] = c286obus[data_w*1 +:data_w];
assign c286ibus[temp_w*2 +:temp_w] = v559obus[temp_w*1 +:temp_w];
assign v559ibus[data_w*1 +:data_w] = c286obus[data_w*2 +:data_w];
assign c286ibus[temp_w*3 +:temp_w] = v703obus[temp_w*1 +:temp_w];
assign v703ibus[data_w*1 +:data_w] = c286obus[data_w*3 +:data_w];
assign c286ibus[temp_w*4 +:temp_w] = v1150obus[temp_w*1 +:temp_w];
assign v1150ibus[data_w*1 +:data_w] = c286obus[data_w*4 +:data_w];
assign c286ibus[temp_w*5 +:temp_w] = v1438obus[temp_w*1 +:temp_w];
assign v1438ibus[data_w*1 +:data_w] = c286obus[data_w*5 +:data_w];
assign c286ibus[temp_w*6 +:temp_w] = v1534obus[temp_w*0 +:temp_w];
assign v1534ibus[data_w*0 +:data_w] = c286obus[data_w*6 +:data_w];
assign c287ibus[temp_w*0 +:temp_w] = v311obus[temp_w*0 +:temp_w];
assign v311ibus[data_w*0 +:data_w] = c287obus[data_w*0 +:data_w];
assign c287ibus[temp_w*1 +:temp_w] = v405obus[temp_w*0 +:temp_w];
assign v405ibus[data_w*0 +:data_w] = c287obus[data_w*1 +:data_w];
assign c287ibus[temp_w*2 +:temp_w] = v560obus[temp_w*1 +:temp_w];
assign v560ibus[data_w*1 +:data_w] = c287obus[data_w*2 +:data_w];
assign c287ibus[temp_w*3 +:temp_w] = v704obus[temp_w*1 +:temp_w];
assign v704ibus[data_w*1 +:data_w] = c287obus[data_w*3 +:data_w];
assign c287ibus[temp_w*4 +:temp_w] = v1151obus[temp_w*1 +:temp_w];
assign v1151ibus[data_w*1 +:data_w] = c287obus[data_w*4 +:data_w];
assign c287ibus[temp_w*5 +:temp_w] = v1439obus[temp_w*1 +:temp_w];
assign v1439ibus[data_w*1 +:data_w] = c287obus[data_w*5 +:data_w];
assign c287ibus[temp_w*6 +:temp_w] = v1535obus[temp_w*0 +:temp_w];
assign v1535ibus[data_w*0 +:data_w] = c287obus[data_w*6 +:data_w];
assign c288ibus[temp_w*0 +:temp_w] = v61obus[temp_w*0 +:temp_w];
assign v61ibus[data_w*0 +:data_w] = c288obus[data_w*0 +:data_w];
assign c288ibus[temp_w*1 +:temp_w] = v239obus[temp_w*1 +:temp_w];
assign v239ibus[data_w*1 +:data_w] = c288obus[data_w*1 +:data_w];
assign c288ibus[temp_w*2 +:temp_w] = v833obus[temp_w*1 +:temp_w];
assign v833ibus[data_w*1 +:data_w] = c288obus[data_w*2 +:data_w];
assign c288ibus[temp_w*3 +:temp_w] = v889obus[temp_w*1 +:temp_w];
assign v889ibus[data_w*1 +:data_w] = c288obus[data_w*3 +:data_w];
assign c288ibus[temp_w*4 +:temp_w] = v1440obus[temp_w*1 +:temp_w];
assign v1440ibus[data_w*1 +:data_w] = c288obus[data_w*4 +:data_w];
assign c288ibus[temp_w*5 +:temp_w] = v1536obus[temp_w*0 +:temp_w];
assign v1536ibus[data_w*0 +:data_w] = c288obus[data_w*5 +:data_w];
assign c289ibus[temp_w*0 +:temp_w] = v62obus[temp_w*0 +:temp_w];
assign v62ibus[data_w*0 +:data_w] = c289obus[data_w*0 +:data_w];
assign c289ibus[temp_w*1 +:temp_w] = v240obus[temp_w*1 +:temp_w];
assign v240ibus[data_w*1 +:data_w] = c289obus[data_w*1 +:data_w];
assign c289ibus[temp_w*2 +:temp_w] = v834obus[temp_w*1 +:temp_w];
assign v834ibus[data_w*1 +:data_w] = c289obus[data_w*2 +:data_w];
assign c289ibus[temp_w*3 +:temp_w] = v890obus[temp_w*1 +:temp_w];
assign v890ibus[data_w*1 +:data_w] = c289obus[data_w*3 +:data_w];
assign c289ibus[temp_w*4 +:temp_w] = v1441obus[temp_w*1 +:temp_w];
assign v1441ibus[data_w*1 +:data_w] = c289obus[data_w*4 +:data_w];
assign c289ibus[temp_w*5 +:temp_w] = v1537obus[temp_w*0 +:temp_w];
assign v1537ibus[data_w*0 +:data_w] = c289obus[data_w*5 +:data_w];
assign c290ibus[temp_w*0 +:temp_w] = v63obus[temp_w*0 +:temp_w];
assign v63ibus[data_w*0 +:data_w] = c290obus[data_w*0 +:data_w];
assign c290ibus[temp_w*1 +:temp_w] = v241obus[temp_w*1 +:temp_w];
assign v241ibus[data_w*1 +:data_w] = c290obus[data_w*1 +:data_w];
assign c290ibus[temp_w*2 +:temp_w] = v835obus[temp_w*1 +:temp_w];
assign v835ibus[data_w*1 +:data_w] = c290obus[data_w*2 +:data_w];
assign c290ibus[temp_w*3 +:temp_w] = v891obus[temp_w*1 +:temp_w];
assign v891ibus[data_w*1 +:data_w] = c290obus[data_w*3 +:data_w];
assign c290ibus[temp_w*4 +:temp_w] = v1442obus[temp_w*1 +:temp_w];
assign v1442ibus[data_w*1 +:data_w] = c290obus[data_w*4 +:data_w];
assign c290ibus[temp_w*5 +:temp_w] = v1538obus[temp_w*0 +:temp_w];
assign v1538ibus[data_w*0 +:data_w] = c290obus[data_w*5 +:data_w];
assign c291ibus[temp_w*0 +:temp_w] = v64obus[temp_w*0 +:temp_w];
assign v64ibus[data_w*0 +:data_w] = c291obus[data_w*0 +:data_w];
assign c291ibus[temp_w*1 +:temp_w] = v242obus[temp_w*1 +:temp_w];
assign v242ibus[data_w*1 +:data_w] = c291obus[data_w*1 +:data_w];
assign c291ibus[temp_w*2 +:temp_w] = v836obus[temp_w*1 +:temp_w];
assign v836ibus[data_w*1 +:data_w] = c291obus[data_w*2 +:data_w];
assign c291ibus[temp_w*3 +:temp_w] = v892obus[temp_w*1 +:temp_w];
assign v892ibus[data_w*1 +:data_w] = c291obus[data_w*3 +:data_w];
assign c291ibus[temp_w*4 +:temp_w] = v1443obus[temp_w*1 +:temp_w];
assign v1443ibus[data_w*1 +:data_w] = c291obus[data_w*4 +:data_w];
assign c291ibus[temp_w*5 +:temp_w] = v1539obus[temp_w*0 +:temp_w];
assign v1539ibus[data_w*0 +:data_w] = c291obus[data_w*5 +:data_w];
assign c292ibus[temp_w*0 +:temp_w] = v65obus[temp_w*0 +:temp_w];
assign v65ibus[data_w*0 +:data_w] = c292obus[data_w*0 +:data_w];
assign c292ibus[temp_w*1 +:temp_w] = v243obus[temp_w*1 +:temp_w];
assign v243ibus[data_w*1 +:data_w] = c292obus[data_w*1 +:data_w];
assign c292ibus[temp_w*2 +:temp_w] = v837obus[temp_w*1 +:temp_w];
assign v837ibus[data_w*1 +:data_w] = c292obus[data_w*2 +:data_w];
assign c292ibus[temp_w*3 +:temp_w] = v893obus[temp_w*1 +:temp_w];
assign v893ibus[data_w*1 +:data_w] = c292obus[data_w*3 +:data_w];
assign c292ibus[temp_w*4 +:temp_w] = v1444obus[temp_w*1 +:temp_w];
assign v1444ibus[data_w*1 +:data_w] = c292obus[data_w*4 +:data_w];
assign c292ibus[temp_w*5 +:temp_w] = v1540obus[temp_w*0 +:temp_w];
assign v1540ibus[data_w*0 +:data_w] = c292obus[data_w*5 +:data_w];
assign c293ibus[temp_w*0 +:temp_w] = v66obus[temp_w*0 +:temp_w];
assign v66ibus[data_w*0 +:data_w] = c293obus[data_w*0 +:data_w];
assign c293ibus[temp_w*1 +:temp_w] = v244obus[temp_w*1 +:temp_w];
assign v244ibus[data_w*1 +:data_w] = c293obus[data_w*1 +:data_w];
assign c293ibus[temp_w*2 +:temp_w] = v838obus[temp_w*1 +:temp_w];
assign v838ibus[data_w*1 +:data_w] = c293obus[data_w*2 +:data_w];
assign c293ibus[temp_w*3 +:temp_w] = v894obus[temp_w*1 +:temp_w];
assign v894ibus[data_w*1 +:data_w] = c293obus[data_w*3 +:data_w];
assign c293ibus[temp_w*4 +:temp_w] = v1445obus[temp_w*1 +:temp_w];
assign v1445ibus[data_w*1 +:data_w] = c293obus[data_w*4 +:data_w];
assign c293ibus[temp_w*5 +:temp_w] = v1541obus[temp_w*0 +:temp_w];
assign v1541ibus[data_w*0 +:data_w] = c293obus[data_w*5 +:data_w];
assign c294ibus[temp_w*0 +:temp_w] = v67obus[temp_w*0 +:temp_w];
assign v67ibus[data_w*0 +:data_w] = c294obus[data_w*0 +:data_w];
assign c294ibus[temp_w*1 +:temp_w] = v245obus[temp_w*1 +:temp_w];
assign v245ibus[data_w*1 +:data_w] = c294obus[data_w*1 +:data_w];
assign c294ibus[temp_w*2 +:temp_w] = v839obus[temp_w*1 +:temp_w];
assign v839ibus[data_w*1 +:data_w] = c294obus[data_w*2 +:data_w];
assign c294ibus[temp_w*3 +:temp_w] = v895obus[temp_w*1 +:temp_w];
assign v895ibus[data_w*1 +:data_w] = c294obus[data_w*3 +:data_w];
assign c294ibus[temp_w*4 +:temp_w] = v1446obus[temp_w*1 +:temp_w];
assign v1446ibus[data_w*1 +:data_w] = c294obus[data_w*4 +:data_w];
assign c294ibus[temp_w*5 +:temp_w] = v1542obus[temp_w*0 +:temp_w];
assign v1542ibus[data_w*0 +:data_w] = c294obus[data_w*5 +:data_w];
assign c295ibus[temp_w*0 +:temp_w] = v68obus[temp_w*0 +:temp_w];
assign v68ibus[data_w*0 +:data_w] = c295obus[data_w*0 +:data_w];
assign c295ibus[temp_w*1 +:temp_w] = v246obus[temp_w*1 +:temp_w];
assign v246ibus[data_w*1 +:data_w] = c295obus[data_w*1 +:data_w];
assign c295ibus[temp_w*2 +:temp_w] = v840obus[temp_w*1 +:temp_w];
assign v840ibus[data_w*1 +:data_w] = c295obus[data_w*2 +:data_w];
assign c295ibus[temp_w*3 +:temp_w] = v896obus[temp_w*1 +:temp_w];
assign v896ibus[data_w*1 +:data_w] = c295obus[data_w*3 +:data_w];
assign c295ibus[temp_w*4 +:temp_w] = v1447obus[temp_w*1 +:temp_w];
assign v1447ibus[data_w*1 +:data_w] = c295obus[data_w*4 +:data_w];
assign c295ibus[temp_w*5 +:temp_w] = v1543obus[temp_w*0 +:temp_w];
assign v1543ibus[data_w*0 +:data_w] = c295obus[data_w*5 +:data_w];
assign c296ibus[temp_w*0 +:temp_w] = v69obus[temp_w*0 +:temp_w];
assign v69ibus[data_w*0 +:data_w] = c296obus[data_w*0 +:data_w];
assign c296ibus[temp_w*1 +:temp_w] = v247obus[temp_w*1 +:temp_w];
assign v247ibus[data_w*1 +:data_w] = c296obus[data_w*1 +:data_w];
assign c296ibus[temp_w*2 +:temp_w] = v841obus[temp_w*1 +:temp_w];
assign v841ibus[data_w*1 +:data_w] = c296obus[data_w*2 +:data_w];
assign c296ibus[temp_w*3 +:temp_w] = v897obus[temp_w*1 +:temp_w];
assign v897ibus[data_w*1 +:data_w] = c296obus[data_w*3 +:data_w];
assign c296ibus[temp_w*4 +:temp_w] = v1448obus[temp_w*1 +:temp_w];
assign v1448ibus[data_w*1 +:data_w] = c296obus[data_w*4 +:data_w];
assign c296ibus[temp_w*5 +:temp_w] = v1544obus[temp_w*0 +:temp_w];
assign v1544ibus[data_w*0 +:data_w] = c296obus[data_w*5 +:data_w];
assign c297ibus[temp_w*0 +:temp_w] = v70obus[temp_w*0 +:temp_w];
assign v70ibus[data_w*0 +:data_w] = c297obus[data_w*0 +:data_w];
assign c297ibus[temp_w*1 +:temp_w] = v248obus[temp_w*1 +:temp_w];
assign v248ibus[data_w*1 +:data_w] = c297obus[data_w*1 +:data_w];
assign c297ibus[temp_w*2 +:temp_w] = v842obus[temp_w*1 +:temp_w];
assign v842ibus[data_w*1 +:data_w] = c297obus[data_w*2 +:data_w];
assign c297ibus[temp_w*3 +:temp_w] = v898obus[temp_w*1 +:temp_w];
assign v898ibus[data_w*1 +:data_w] = c297obus[data_w*3 +:data_w];
assign c297ibus[temp_w*4 +:temp_w] = v1449obus[temp_w*1 +:temp_w];
assign v1449ibus[data_w*1 +:data_w] = c297obus[data_w*4 +:data_w];
assign c297ibus[temp_w*5 +:temp_w] = v1545obus[temp_w*0 +:temp_w];
assign v1545ibus[data_w*0 +:data_w] = c297obus[data_w*5 +:data_w];
assign c298ibus[temp_w*0 +:temp_w] = v71obus[temp_w*0 +:temp_w];
assign v71ibus[data_w*0 +:data_w] = c298obus[data_w*0 +:data_w];
assign c298ibus[temp_w*1 +:temp_w] = v249obus[temp_w*1 +:temp_w];
assign v249ibus[data_w*1 +:data_w] = c298obus[data_w*1 +:data_w];
assign c298ibus[temp_w*2 +:temp_w] = v843obus[temp_w*1 +:temp_w];
assign v843ibus[data_w*1 +:data_w] = c298obus[data_w*2 +:data_w];
assign c298ibus[temp_w*3 +:temp_w] = v899obus[temp_w*1 +:temp_w];
assign v899ibus[data_w*1 +:data_w] = c298obus[data_w*3 +:data_w];
assign c298ibus[temp_w*4 +:temp_w] = v1450obus[temp_w*1 +:temp_w];
assign v1450ibus[data_w*1 +:data_w] = c298obus[data_w*4 +:data_w];
assign c298ibus[temp_w*5 +:temp_w] = v1546obus[temp_w*0 +:temp_w];
assign v1546ibus[data_w*0 +:data_w] = c298obus[data_w*5 +:data_w];
assign c299ibus[temp_w*0 +:temp_w] = v72obus[temp_w*0 +:temp_w];
assign v72ibus[data_w*0 +:data_w] = c299obus[data_w*0 +:data_w];
assign c299ibus[temp_w*1 +:temp_w] = v250obus[temp_w*1 +:temp_w];
assign v250ibus[data_w*1 +:data_w] = c299obus[data_w*1 +:data_w];
assign c299ibus[temp_w*2 +:temp_w] = v844obus[temp_w*1 +:temp_w];
assign v844ibus[data_w*1 +:data_w] = c299obus[data_w*2 +:data_w];
assign c299ibus[temp_w*3 +:temp_w] = v900obus[temp_w*1 +:temp_w];
assign v900ibus[data_w*1 +:data_w] = c299obus[data_w*3 +:data_w];
assign c299ibus[temp_w*4 +:temp_w] = v1451obus[temp_w*1 +:temp_w];
assign v1451ibus[data_w*1 +:data_w] = c299obus[data_w*4 +:data_w];
assign c299ibus[temp_w*5 +:temp_w] = v1547obus[temp_w*0 +:temp_w];
assign v1547ibus[data_w*0 +:data_w] = c299obus[data_w*5 +:data_w];
assign c300ibus[temp_w*0 +:temp_w] = v73obus[temp_w*0 +:temp_w];
assign v73ibus[data_w*0 +:data_w] = c300obus[data_w*0 +:data_w];
assign c300ibus[temp_w*1 +:temp_w] = v251obus[temp_w*1 +:temp_w];
assign v251ibus[data_w*1 +:data_w] = c300obus[data_w*1 +:data_w];
assign c300ibus[temp_w*2 +:temp_w] = v845obus[temp_w*1 +:temp_w];
assign v845ibus[data_w*1 +:data_w] = c300obus[data_w*2 +:data_w];
assign c300ibus[temp_w*3 +:temp_w] = v901obus[temp_w*1 +:temp_w];
assign v901ibus[data_w*1 +:data_w] = c300obus[data_w*3 +:data_w];
assign c300ibus[temp_w*4 +:temp_w] = v1452obus[temp_w*1 +:temp_w];
assign v1452ibus[data_w*1 +:data_w] = c300obus[data_w*4 +:data_w];
assign c300ibus[temp_w*5 +:temp_w] = v1548obus[temp_w*0 +:temp_w];
assign v1548ibus[data_w*0 +:data_w] = c300obus[data_w*5 +:data_w];
assign c301ibus[temp_w*0 +:temp_w] = v74obus[temp_w*0 +:temp_w];
assign v74ibus[data_w*0 +:data_w] = c301obus[data_w*0 +:data_w];
assign c301ibus[temp_w*1 +:temp_w] = v252obus[temp_w*1 +:temp_w];
assign v252ibus[data_w*1 +:data_w] = c301obus[data_w*1 +:data_w];
assign c301ibus[temp_w*2 +:temp_w] = v846obus[temp_w*1 +:temp_w];
assign v846ibus[data_w*1 +:data_w] = c301obus[data_w*2 +:data_w];
assign c301ibus[temp_w*3 +:temp_w] = v902obus[temp_w*1 +:temp_w];
assign v902ibus[data_w*1 +:data_w] = c301obus[data_w*3 +:data_w];
assign c301ibus[temp_w*4 +:temp_w] = v1453obus[temp_w*1 +:temp_w];
assign v1453ibus[data_w*1 +:data_w] = c301obus[data_w*4 +:data_w];
assign c301ibus[temp_w*5 +:temp_w] = v1549obus[temp_w*0 +:temp_w];
assign v1549ibus[data_w*0 +:data_w] = c301obus[data_w*5 +:data_w];
assign c302ibus[temp_w*0 +:temp_w] = v75obus[temp_w*0 +:temp_w];
assign v75ibus[data_w*0 +:data_w] = c302obus[data_w*0 +:data_w];
assign c302ibus[temp_w*1 +:temp_w] = v253obus[temp_w*1 +:temp_w];
assign v253ibus[data_w*1 +:data_w] = c302obus[data_w*1 +:data_w];
assign c302ibus[temp_w*2 +:temp_w] = v847obus[temp_w*1 +:temp_w];
assign v847ibus[data_w*1 +:data_w] = c302obus[data_w*2 +:data_w];
assign c302ibus[temp_w*3 +:temp_w] = v903obus[temp_w*1 +:temp_w];
assign v903ibus[data_w*1 +:data_w] = c302obus[data_w*3 +:data_w];
assign c302ibus[temp_w*4 +:temp_w] = v1454obus[temp_w*1 +:temp_w];
assign v1454ibus[data_w*1 +:data_w] = c302obus[data_w*4 +:data_w];
assign c302ibus[temp_w*5 +:temp_w] = v1550obus[temp_w*0 +:temp_w];
assign v1550ibus[data_w*0 +:data_w] = c302obus[data_w*5 +:data_w];
assign c303ibus[temp_w*0 +:temp_w] = v76obus[temp_w*0 +:temp_w];
assign v76ibus[data_w*0 +:data_w] = c303obus[data_w*0 +:data_w];
assign c303ibus[temp_w*1 +:temp_w] = v254obus[temp_w*1 +:temp_w];
assign v254ibus[data_w*1 +:data_w] = c303obus[data_w*1 +:data_w];
assign c303ibus[temp_w*2 +:temp_w] = v848obus[temp_w*1 +:temp_w];
assign v848ibus[data_w*1 +:data_w] = c303obus[data_w*2 +:data_w];
assign c303ibus[temp_w*3 +:temp_w] = v904obus[temp_w*1 +:temp_w];
assign v904ibus[data_w*1 +:data_w] = c303obus[data_w*3 +:data_w];
assign c303ibus[temp_w*4 +:temp_w] = v1455obus[temp_w*1 +:temp_w];
assign v1455ibus[data_w*1 +:data_w] = c303obus[data_w*4 +:data_w];
assign c303ibus[temp_w*5 +:temp_w] = v1551obus[temp_w*0 +:temp_w];
assign v1551ibus[data_w*0 +:data_w] = c303obus[data_w*5 +:data_w];
assign c304ibus[temp_w*0 +:temp_w] = v77obus[temp_w*0 +:temp_w];
assign v77ibus[data_w*0 +:data_w] = c304obus[data_w*0 +:data_w];
assign c304ibus[temp_w*1 +:temp_w] = v255obus[temp_w*1 +:temp_w];
assign v255ibus[data_w*1 +:data_w] = c304obus[data_w*1 +:data_w];
assign c304ibus[temp_w*2 +:temp_w] = v849obus[temp_w*1 +:temp_w];
assign v849ibus[data_w*1 +:data_w] = c304obus[data_w*2 +:data_w];
assign c304ibus[temp_w*3 +:temp_w] = v905obus[temp_w*1 +:temp_w];
assign v905ibus[data_w*1 +:data_w] = c304obus[data_w*3 +:data_w];
assign c304ibus[temp_w*4 +:temp_w] = v1456obus[temp_w*1 +:temp_w];
assign v1456ibus[data_w*1 +:data_w] = c304obus[data_w*4 +:data_w];
assign c304ibus[temp_w*5 +:temp_w] = v1552obus[temp_w*0 +:temp_w];
assign v1552ibus[data_w*0 +:data_w] = c304obus[data_w*5 +:data_w];
assign c305ibus[temp_w*0 +:temp_w] = v78obus[temp_w*0 +:temp_w];
assign v78ibus[data_w*0 +:data_w] = c305obus[data_w*0 +:data_w];
assign c305ibus[temp_w*1 +:temp_w] = v256obus[temp_w*1 +:temp_w];
assign v256ibus[data_w*1 +:data_w] = c305obus[data_w*1 +:data_w];
assign c305ibus[temp_w*2 +:temp_w] = v850obus[temp_w*1 +:temp_w];
assign v850ibus[data_w*1 +:data_w] = c305obus[data_w*2 +:data_w];
assign c305ibus[temp_w*3 +:temp_w] = v906obus[temp_w*1 +:temp_w];
assign v906ibus[data_w*1 +:data_w] = c305obus[data_w*3 +:data_w];
assign c305ibus[temp_w*4 +:temp_w] = v1457obus[temp_w*1 +:temp_w];
assign v1457ibus[data_w*1 +:data_w] = c305obus[data_w*4 +:data_w];
assign c305ibus[temp_w*5 +:temp_w] = v1553obus[temp_w*0 +:temp_w];
assign v1553ibus[data_w*0 +:data_w] = c305obus[data_w*5 +:data_w];
assign c306ibus[temp_w*0 +:temp_w] = v79obus[temp_w*0 +:temp_w];
assign v79ibus[data_w*0 +:data_w] = c306obus[data_w*0 +:data_w];
assign c306ibus[temp_w*1 +:temp_w] = v257obus[temp_w*1 +:temp_w];
assign v257ibus[data_w*1 +:data_w] = c306obus[data_w*1 +:data_w];
assign c306ibus[temp_w*2 +:temp_w] = v851obus[temp_w*1 +:temp_w];
assign v851ibus[data_w*1 +:data_w] = c306obus[data_w*2 +:data_w];
assign c306ibus[temp_w*3 +:temp_w] = v907obus[temp_w*1 +:temp_w];
assign v907ibus[data_w*1 +:data_w] = c306obus[data_w*3 +:data_w];
assign c306ibus[temp_w*4 +:temp_w] = v1458obus[temp_w*1 +:temp_w];
assign v1458ibus[data_w*1 +:data_w] = c306obus[data_w*4 +:data_w];
assign c306ibus[temp_w*5 +:temp_w] = v1554obus[temp_w*0 +:temp_w];
assign v1554ibus[data_w*0 +:data_w] = c306obus[data_w*5 +:data_w];
assign c307ibus[temp_w*0 +:temp_w] = v80obus[temp_w*0 +:temp_w];
assign v80ibus[data_w*0 +:data_w] = c307obus[data_w*0 +:data_w];
assign c307ibus[temp_w*1 +:temp_w] = v258obus[temp_w*1 +:temp_w];
assign v258ibus[data_w*1 +:data_w] = c307obus[data_w*1 +:data_w];
assign c307ibus[temp_w*2 +:temp_w] = v852obus[temp_w*1 +:temp_w];
assign v852ibus[data_w*1 +:data_w] = c307obus[data_w*2 +:data_w];
assign c307ibus[temp_w*3 +:temp_w] = v908obus[temp_w*1 +:temp_w];
assign v908ibus[data_w*1 +:data_w] = c307obus[data_w*3 +:data_w];
assign c307ibus[temp_w*4 +:temp_w] = v1459obus[temp_w*1 +:temp_w];
assign v1459ibus[data_w*1 +:data_w] = c307obus[data_w*4 +:data_w];
assign c307ibus[temp_w*5 +:temp_w] = v1555obus[temp_w*0 +:temp_w];
assign v1555ibus[data_w*0 +:data_w] = c307obus[data_w*5 +:data_w];
assign c308ibus[temp_w*0 +:temp_w] = v81obus[temp_w*0 +:temp_w];
assign v81ibus[data_w*0 +:data_w] = c308obus[data_w*0 +:data_w];
assign c308ibus[temp_w*1 +:temp_w] = v259obus[temp_w*1 +:temp_w];
assign v259ibus[data_w*1 +:data_w] = c308obus[data_w*1 +:data_w];
assign c308ibus[temp_w*2 +:temp_w] = v853obus[temp_w*1 +:temp_w];
assign v853ibus[data_w*1 +:data_w] = c308obus[data_w*2 +:data_w];
assign c308ibus[temp_w*3 +:temp_w] = v909obus[temp_w*1 +:temp_w];
assign v909ibus[data_w*1 +:data_w] = c308obus[data_w*3 +:data_w];
assign c308ibus[temp_w*4 +:temp_w] = v1460obus[temp_w*1 +:temp_w];
assign v1460ibus[data_w*1 +:data_w] = c308obus[data_w*4 +:data_w];
assign c308ibus[temp_w*5 +:temp_w] = v1556obus[temp_w*0 +:temp_w];
assign v1556ibus[data_w*0 +:data_w] = c308obus[data_w*5 +:data_w];
assign c309ibus[temp_w*0 +:temp_w] = v82obus[temp_w*0 +:temp_w];
assign v82ibus[data_w*0 +:data_w] = c309obus[data_w*0 +:data_w];
assign c309ibus[temp_w*1 +:temp_w] = v260obus[temp_w*1 +:temp_w];
assign v260ibus[data_w*1 +:data_w] = c309obus[data_w*1 +:data_w];
assign c309ibus[temp_w*2 +:temp_w] = v854obus[temp_w*1 +:temp_w];
assign v854ibus[data_w*1 +:data_w] = c309obus[data_w*2 +:data_w];
assign c309ibus[temp_w*3 +:temp_w] = v910obus[temp_w*1 +:temp_w];
assign v910ibus[data_w*1 +:data_w] = c309obus[data_w*3 +:data_w];
assign c309ibus[temp_w*4 +:temp_w] = v1461obus[temp_w*1 +:temp_w];
assign v1461ibus[data_w*1 +:data_w] = c309obus[data_w*4 +:data_w];
assign c309ibus[temp_w*5 +:temp_w] = v1557obus[temp_w*0 +:temp_w];
assign v1557ibus[data_w*0 +:data_w] = c309obus[data_w*5 +:data_w];
assign c310ibus[temp_w*0 +:temp_w] = v83obus[temp_w*0 +:temp_w];
assign v83ibus[data_w*0 +:data_w] = c310obus[data_w*0 +:data_w];
assign c310ibus[temp_w*1 +:temp_w] = v261obus[temp_w*1 +:temp_w];
assign v261ibus[data_w*1 +:data_w] = c310obus[data_w*1 +:data_w];
assign c310ibus[temp_w*2 +:temp_w] = v855obus[temp_w*1 +:temp_w];
assign v855ibus[data_w*1 +:data_w] = c310obus[data_w*2 +:data_w];
assign c310ibus[temp_w*3 +:temp_w] = v911obus[temp_w*1 +:temp_w];
assign v911ibus[data_w*1 +:data_w] = c310obus[data_w*3 +:data_w];
assign c310ibus[temp_w*4 +:temp_w] = v1462obus[temp_w*1 +:temp_w];
assign v1462ibus[data_w*1 +:data_w] = c310obus[data_w*4 +:data_w];
assign c310ibus[temp_w*5 +:temp_w] = v1558obus[temp_w*0 +:temp_w];
assign v1558ibus[data_w*0 +:data_w] = c310obus[data_w*5 +:data_w];
assign c311ibus[temp_w*0 +:temp_w] = v84obus[temp_w*0 +:temp_w];
assign v84ibus[data_w*0 +:data_w] = c311obus[data_w*0 +:data_w];
assign c311ibus[temp_w*1 +:temp_w] = v262obus[temp_w*1 +:temp_w];
assign v262ibus[data_w*1 +:data_w] = c311obus[data_w*1 +:data_w];
assign c311ibus[temp_w*2 +:temp_w] = v856obus[temp_w*1 +:temp_w];
assign v856ibus[data_w*1 +:data_w] = c311obus[data_w*2 +:data_w];
assign c311ibus[temp_w*3 +:temp_w] = v912obus[temp_w*1 +:temp_w];
assign v912ibus[data_w*1 +:data_w] = c311obus[data_w*3 +:data_w];
assign c311ibus[temp_w*4 +:temp_w] = v1463obus[temp_w*1 +:temp_w];
assign v1463ibus[data_w*1 +:data_w] = c311obus[data_w*4 +:data_w];
assign c311ibus[temp_w*5 +:temp_w] = v1559obus[temp_w*0 +:temp_w];
assign v1559ibus[data_w*0 +:data_w] = c311obus[data_w*5 +:data_w];
assign c312ibus[temp_w*0 +:temp_w] = v85obus[temp_w*0 +:temp_w];
assign v85ibus[data_w*0 +:data_w] = c312obus[data_w*0 +:data_w];
assign c312ibus[temp_w*1 +:temp_w] = v263obus[temp_w*1 +:temp_w];
assign v263ibus[data_w*1 +:data_w] = c312obus[data_w*1 +:data_w];
assign c312ibus[temp_w*2 +:temp_w] = v857obus[temp_w*1 +:temp_w];
assign v857ibus[data_w*1 +:data_w] = c312obus[data_w*2 +:data_w];
assign c312ibus[temp_w*3 +:temp_w] = v913obus[temp_w*1 +:temp_w];
assign v913ibus[data_w*1 +:data_w] = c312obus[data_w*3 +:data_w];
assign c312ibus[temp_w*4 +:temp_w] = v1464obus[temp_w*1 +:temp_w];
assign v1464ibus[data_w*1 +:data_w] = c312obus[data_w*4 +:data_w];
assign c312ibus[temp_w*5 +:temp_w] = v1560obus[temp_w*0 +:temp_w];
assign v1560ibus[data_w*0 +:data_w] = c312obus[data_w*5 +:data_w];
assign c313ibus[temp_w*0 +:temp_w] = v86obus[temp_w*0 +:temp_w];
assign v86ibus[data_w*0 +:data_w] = c313obus[data_w*0 +:data_w];
assign c313ibus[temp_w*1 +:temp_w] = v264obus[temp_w*1 +:temp_w];
assign v264ibus[data_w*1 +:data_w] = c313obus[data_w*1 +:data_w];
assign c313ibus[temp_w*2 +:temp_w] = v858obus[temp_w*1 +:temp_w];
assign v858ibus[data_w*1 +:data_w] = c313obus[data_w*2 +:data_w];
assign c313ibus[temp_w*3 +:temp_w] = v914obus[temp_w*1 +:temp_w];
assign v914ibus[data_w*1 +:data_w] = c313obus[data_w*3 +:data_w];
assign c313ibus[temp_w*4 +:temp_w] = v1465obus[temp_w*1 +:temp_w];
assign v1465ibus[data_w*1 +:data_w] = c313obus[data_w*4 +:data_w];
assign c313ibus[temp_w*5 +:temp_w] = v1561obus[temp_w*0 +:temp_w];
assign v1561ibus[data_w*0 +:data_w] = c313obus[data_w*5 +:data_w];
assign c314ibus[temp_w*0 +:temp_w] = v87obus[temp_w*0 +:temp_w];
assign v87ibus[data_w*0 +:data_w] = c314obus[data_w*0 +:data_w];
assign c314ibus[temp_w*1 +:temp_w] = v265obus[temp_w*1 +:temp_w];
assign v265ibus[data_w*1 +:data_w] = c314obus[data_w*1 +:data_w];
assign c314ibus[temp_w*2 +:temp_w] = v859obus[temp_w*1 +:temp_w];
assign v859ibus[data_w*1 +:data_w] = c314obus[data_w*2 +:data_w];
assign c314ibus[temp_w*3 +:temp_w] = v915obus[temp_w*1 +:temp_w];
assign v915ibus[data_w*1 +:data_w] = c314obus[data_w*3 +:data_w];
assign c314ibus[temp_w*4 +:temp_w] = v1466obus[temp_w*1 +:temp_w];
assign v1466ibus[data_w*1 +:data_w] = c314obus[data_w*4 +:data_w];
assign c314ibus[temp_w*5 +:temp_w] = v1562obus[temp_w*0 +:temp_w];
assign v1562ibus[data_w*0 +:data_w] = c314obus[data_w*5 +:data_w];
assign c315ibus[temp_w*0 +:temp_w] = v88obus[temp_w*0 +:temp_w];
assign v88ibus[data_w*0 +:data_w] = c315obus[data_w*0 +:data_w];
assign c315ibus[temp_w*1 +:temp_w] = v266obus[temp_w*1 +:temp_w];
assign v266ibus[data_w*1 +:data_w] = c315obus[data_w*1 +:data_w];
assign c315ibus[temp_w*2 +:temp_w] = v860obus[temp_w*1 +:temp_w];
assign v860ibus[data_w*1 +:data_w] = c315obus[data_w*2 +:data_w];
assign c315ibus[temp_w*3 +:temp_w] = v916obus[temp_w*1 +:temp_w];
assign v916ibus[data_w*1 +:data_w] = c315obus[data_w*3 +:data_w];
assign c315ibus[temp_w*4 +:temp_w] = v1467obus[temp_w*1 +:temp_w];
assign v1467ibus[data_w*1 +:data_w] = c315obus[data_w*4 +:data_w];
assign c315ibus[temp_w*5 +:temp_w] = v1563obus[temp_w*0 +:temp_w];
assign v1563ibus[data_w*0 +:data_w] = c315obus[data_w*5 +:data_w];
assign c316ibus[temp_w*0 +:temp_w] = v89obus[temp_w*0 +:temp_w];
assign v89ibus[data_w*0 +:data_w] = c316obus[data_w*0 +:data_w];
assign c316ibus[temp_w*1 +:temp_w] = v267obus[temp_w*1 +:temp_w];
assign v267ibus[data_w*1 +:data_w] = c316obus[data_w*1 +:data_w];
assign c316ibus[temp_w*2 +:temp_w] = v861obus[temp_w*1 +:temp_w];
assign v861ibus[data_w*1 +:data_w] = c316obus[data_w*2 +:data_w];
assign c316ibus[temp_w*3 +:temp_w] = v917obus[temp_w*1 +:temp_w];
assign v917ibus[data_w*1 +:data_w] = c316obus[data_w*3 +:data_w];
assign c316ibus[temp_w*4 +:temp_w] = v1468obus[temp_w*1 +:temp_w];
assign v1468ibus[data_w*1 +:data_w] = c316obus[data_w*4 +:data_w];
assign c316ibus[temp_w*5 +:temp_w] = v1564obus[temp_w*0 +:temp_w];
assign v1564ibus[data_w*0 +:data_w] = c316obus[data_w*5 +:data_w];
assign c317ibus[temp_w*0 +:temp_w] = v90obus[temp_w*0 +:temp_w];
assign v90ibus[data_w*0 +:data_w] = c317obus[data_w*0 +:data_w];
assign c317ibus[temp_w*1 +:temp_w] = v268obus[temp_w*1 +:temp_w];
assign v268ibus[data_w*1 +:data_w] = c317obus[data_w*1 +:data_w];
assign c317ibus[temp_w*2 +:temp_w] = v862obus[temp_w*1 +:temp_w];
assign v862ibus[data_w*1 +:data_w] = c317obus[data_w*2 +:data_w];
assign c317ibus[temp_w*3 +:temp_w] = v918obus[temp_w*1 +:temp_w];
assign v918ibus[data_w*1 +:data_w] = c317obus[data_w*3 +:data_w];
assign c317ibus[temp_w*4 +:temp_w] = v1469obus[temp_w*1 +:temp_w];
assign v1469ibus[data_w*1 +:data_w] = c317obus[data_w*4 +:data_w];
assign c317ibus[temp_w*5 +:temp_w] = v1565obus[temp_w*0 +:temp_w];
assign v1565ibus[data_w*0 +:data_w] = c317obus[data_w*5 +:data_w];
assign c318ibus[temp_w*0 +:temp_w] = v91obus[temp_w*0 +:temp_w];
assign v91ibus[data_w*0 +:data_w] = c318obus[data_w*0 +:data_w];
assign c318ibus[temp_w*1 +:temp_w] = v269obus[temp_w*1 +:temp_w];
assign v269ibus[data_w*1 +:data_w] = c318obus[data_w*1 +:data_w];
assign c318ibus[temp_w*2 +:temp_w] = v863obus[temp_w*1 +:temp_w];
assign v863ibus[data_w*1 +:data_w] = c318obus[data_w*2 +:data_w];
assign c318ibus[temp_w*3 +:temp_w] = v919obus[temp_w*1 +:temp_w];
assign v919ibus[data_w*1 +:data_w] = c318obus[data_w*3 +:data_w];
assign c318ibus[temp_w*4 +:temp_w] = v1470obus[temp_w*1 +:temp_w];
assign v1470ibus[data_w*1 +:data_w] = c318obus[data_w*4 +:data_w];
assign c318ibus[temp_w*5 +:temp_w] = v1566obus[temp_w*0 +:temp_w];
assign v1566ibus[data_w*0 +:data_w] = c318obus[data_w*5 +:data_w];
assign c319ibus[temp_w*0 +:temp_w] = v92obus[temp_w*0 +:temp_w];
assign v92ibus[data_w*0 +:data_w] = c319obus[data_w*0 +:data_w];
assign c319ibus[temp_w*1 +:temp_w] = v270obus[temp_w*1 +:temp_w];
assign v270ibus[data_w*1 +:data_w] = c319obus[data_w*1 +:data_w];
assign c319ibus[temp_w*2 +:temp_w] = v768obus[temp_w*1 +:temp_w];
assign v768ibus[data_w*1 +:data_w] = c319obus[data_w*2 +:data_w];
assign c319ibus[temp_w*3 +:temp_w] = v920obus[temp_w*1 +:temp_w];
assign v920ibus[data_w*1 +:data_w] = c319obus[data_w*3 +:data_w];
assign c319ibus[temp_w*4 +:temp_w] = v1471obus[temp_w*1 +:temp_w];
assign v1471ibus[data_w*1 +:data_w] = c319obus[data_w*4 +:data_w];
assign c319ibus[temp_w*5 +:temp_w] = v1567obus[temp_w*0 +:temp_w];
assign v1567ibus[data_w*0 +:data_w] = c319obus[data_w*5 +:data_w];
assign c320ibus[temp_w*0 +:temp_w] = v93obus[temp_w*0 +:temp_w];
assign v93ibus[data_w*0 +:data_w] = c320obus[data_w*0 +:data_w];
assign c320ibus[temp_w*1 +:temp_w] = v271obus[temp_w*1 +:temp_w];
assign v271ibus[data_w*1 +:data_w] = c320obus[data_w*1 +:data_w];
assign c320ibus[temp_w*2 +:temp_w] = v769obus[temp_w*1 +:temp_w];
assign v769ibus[data_w*1 +:data_w] = c320obus[data_w*2 +:data_w];
assign c320ibus[temp_w*3 +:temp_w] = v921obus[temp_w*1 +:temp_w];
assign v921ibus[data_w*1 +:data_w] = c320obus[data_w*3 +:data_w];
assign c320ibus[temp_w*4 +:temp_w] = v1472obus[temp_w*1 +:temp_w];
assign v1472ibus[data_w*1 +:data_w] = c320obus[data_w*4 +:data_w];
assign c320ibus[temp_w*5 +:temp_w] = v1568obus[temp_w*0 +:temp_w];
assign v1568ibus[data_w*0 +:data_w] = c320obus[data_w*5 +:data_w];
assign c321ibus[temp_w*0 +:temp_w] = v94obus[temp_w*0 +:temp_w];
assign v94ibus[data_w*0 +:data_w] = c321obus[data_w*0 +:data_w];
assign c321ibus[temp_w*1 +:temp_w] = v272obus[temp_w*1 +:temp_w];
assign v272ibus[data_w*1 +:data_w] = c321obus[data_w*1 +:data_w];
assign c321ibus[temp_w*2 +:temp_w] = v770obus[temp_w*1 +:temp_w];
assign v770ibus[data_w*1 +:data_w] = c321obus[data_w*2 +:data_w];
assign c321ibus[temp_w*3 +:temp_w] = v922obus[temp_w*1 +:temp_w];
assign v922ibus[data_w*1 +:data_w] = c321obus[data_w*3 +:data_w];
assign c321ibus[temp_w*4 +:temp_w] = v1473obus[temp_w*1 +:temp_w];
assign v1473ibus[data_w*1 +:data_w] = c321obus[data_w*4 +:data_w];
assign c321ibus[temp_w*5 +:temp_w] = v1569obus[temp_w*0 +:temp_w];
assign v1569ibus[data_w*0 +:data_w] = c321obus[data_w*5 +:data_w];
assign c322ibus[temp_w*0 +:temp_w] = v95obus[temp_w*0 +:temp_w];
assign v95ibus[data_w*0 +:data_w] = c322obus[data_w*0 +:data_w];
assign c322ibus[temp_w*1 +:temp_w] = v273obus[temp_w*1 +:temp_w];
assign v273ibus[data_w*1 +:data_w] = c322obus[data_w*1 +:data_w];
assign c322ibus[temp_w*2 +:temp_w] = v771obus[temp_w*1 +:temp_w];
assign v771ibus[data_w*1 +:data_w] = c322obus[data_w*2 +:data_w];
assign c322ibus[temp_w*3 +:temp_w] = v923obus[temp_w*1 +:temp_w];
assign v923ibus[data_w*1 +:data_w] = c322obus[data_w*3 +:data_w];
assign c322ibus[temp_w*4 +:temp_w] = v1474obus[temp_w*1 +:temp_w];
assign v1474ibus[data_w*1 +:data_w] = c322obus[data_w*4 +:data_w];
assign c322ibus[temp_w*5 +:temp_w] = v1570obus[temp_w*0 +:temp_w];
assign v1570ibus[data_w*0 +:data_w] = c322obus[data_w*5 +:data_w];
assign c323ibus[temp_w*0 +:temp_w] = v0obus[temp_w*0 +:temp_w];
assign v0ibus[data_w*0 +:data_w] = c323obus[data_w*0 +:data_w];
assign c323ibus[temp_w*1 +:temp_w] = v274obus[temp_w*1 +:temp_w];
assign v274ibus[data_w*1 +:data_w] = c323obus[data_w*1 +:data_w];
assign c323ibus[temp_w*2 +:temp_w] = v772obus[temp_w*1 +:temp_w];
assign v772ibus[data_w*1 +:data_w] = c323obus[data_w*2 +:data_w];
assign c323ibus[temp_w*3 +:temp_w] = v924obus[temp_w*1 +:temp_w];
assign v924ibus[data_w*1 +:data_w] = c323obus[data_w*3 +:data_w];
assign c323ibus[temp_w*4 +:temp_w] = v1475obus[temp_w*1 +:temp_w];
assign v1475ibus[data_w*1 +:data_w] = c323obus[data_w*4 +:data_w];
assign c323ibus[temp_w*5 +:temp_w] = v1571obus[temp_w*0 +:temp_w];
assign v1571ibus[data_w*0 +:data_w] = c323obus[data_w*5 +:data_w];
assign c324ibus[temp_w*0 +:temp_w] = v1obus[temp_w*0 +:temp_w];
assign v1ibus[data_w*0 +:data_w] = c324obus[data_w*0 +:data_w];
assign c324ibus[temp_w*1 +:temp_w] = v275obus[temp_w*1 +:temp_w];
assign v275ibus[data_w*1 +:data_w] = c324obus[data_w*1 +:data_w];
assign c324ibus[temp_w*2 +:temp_w] = v773obus[temp_w*1 +:temp_w];
assign v773ibus[data_w*1 +:data_w] = c324obus[data_w*2 +:data_w];
assign c324ibus[temp_w*3 +:temp_w] = v925obus[temp_w*1 +:temp_w];
assign v925ibus[data_w*1 +:data_w] = c324obus[data_w*3 +:data_w];
assign c324ibus[temp_w*4 +:temp_w] = v1476obus[temp_w*1 +:temp_w];
assign v1476ibus[data_w*1 +:data_w] = c324obus[data_w*4 +:data_w];
assign c324ibus[temp_w*5 +:temp_w] = v1572obus[temp_w*0 +:temp_w];
assign v1572ibus[data_w*0 +:data_w] = c324obus[data_w*5 +:data_w];
assign c325ibus[temp_w*0 +:temp_w] = v2obus[temp_w*0 +:temp_w];
assign v2ibus[data_w*0 +:data_w] = c325obus[data_w*0 +:data_w];
assign c325ibus[temp_w*1 +:temp_w] = v276obus[temp_w*1 +:temp_w];
assign v276ibus[data_w*1 +:data_w] = c325obus[data_w*1 +:data_w];
assign c325ibus[temp_w*2 +:temp_w] = v774obus[temp_w*1 +:temp_w];
assign v774ibus[data_w*1 +:data_w] = c325obus[data_w*2 +:data_w];
assign c325ibus[temp_w*3 +:temp_w] = v926obus[temp_w*1 +:temp_w];
assign v926ibus[data_w*1 +:data_w] = c325obus[data_w*3 +:data_w];
assign c325ibus[temp_w*4 +:temp_w] = v1477obus[temp_w*1 +:temp_w];
assign v1477ibus[data_w*1 +:data_w] = c325obus[data_w*4 +:data_w];
assign c325ibus[temp_w*5 +:temp_w] = v1573obus[temp_w*0 +:temp_w];
assign v1573ibus[data_w*0 +:data_w] = c325obus[data_w*5 +:data_w];
assign c326ibus[temp_w*0 +:temp_w] = v3obus[temp_w*0 +:temp_w];
assign v3ibus[data_w*0 +:data_w] = c326obus[data_w*0 +:data_w];
assign c326ibus[temp_w*1 +:temp_w] = v277obus[temp_w*1 +:temp_w];
assign v277ibus[data_w*1 +:data_w] = c326obus[data_w*1 +:data_w];
assign c326ibus[temp_w*2 +:temp_w] = v775obus[temp_w*1 +:temp_w];
assign v775ibus[data_w*1 +:data_w] = c326obus[data_w*2 +:data_w];
assign c326ibus[temp_w*3 +:temp_w] = v927obus[temp_w*1 +:temp_w];
assign v927ibus[data_w*1 +:data_w] = c326obus[data_w*3 +:data_w];
assign c326ibus[temp_w*4 +:temp_w] = v1478obus[temp_w*1 +:temp_w];
assign v1478ibus[data_w*1 +:data_w] = c326obus[data_w*4 +:data_w];
assign c326ibus[temp_w*5 +:temp_w] = v1574obus[temp_w*0 +:temp_w];
assign v1574ibus[data_w*0 +:data_w] = c326obus[data_w*5 +:data_w];
assign c327ibus[temp_w*0 +:temp_w] = v4obus[temp_w*0 +:temp_w];
assign v4ibus[data_w*0 +:data_w] = c327obus[data_w*0 +:data_w];
assign c327ibus[temp_w*1 +:temp_w] = v278obus[temp_w*1 +:temp_w];
assign v278ibus[data_w*1 +:data_w] = c327obus[data_w*1 +:data_w];
assign c327ibus[temp_w*2 +:temp_w] = v776obus[temp_w*1 +:temp_w];
assign v776ibus[data_w*1 +:data_w] = c327obus[data_w*2 +:data_w];
assign c327ibus[temp_w*3 +:temp_w] = v928obus[temp_w*1 +:temp_w];
assign v928ibus[data_w*1 +:data_w] = c327obus[data_w*3 +:data_w];
assign c327ibus[temp_w*4 +:temp_w] = v1479obus[temp_w*1 +:temp_w];
assign v1479ibus[data_w*1 +:data_w] = c327obus[data_w*4 +:data_w];
assign c327ibus[temp_w*5 +:temp_w] = v1575obus[temp_w*0 +:temp_w];
assign v1575ibus[data_w*0 +:data_w] = c327obus[data_w*5 +:data_w];
assign c328ibus[temp_w*0 +:temp_w] = v5obus[temp_w*0 +:temp_w];
assign v5ibus[data_w*0 +:data_w] = c328obus[data_w*0 +:data_w];
assign c328ibus[temp_w*1 +:temp_w] = v279obus[temp_w*1 +:temp_w];
assign v279ibus[data_w*1 +:data_w] = c328obus[data_w*1 +:data_w];
assign c328ibus[temp_w*2 +:temp_w] = v777obus[temp_w*1 +:temp_w];
assign v777ibus[data_w*1 +:data_w] = c328obus[data_w*2 +:data_w];
assign c328ibus[temp_w*3 +:temp_w] = v929obus[temp_w*1 +:temp_w];
assign v929ibus[data_w*1 +:data_w] = c328obus[data_w*3 +:data_w];
assign c328ibus[temp_w*4 +:temp_w] = v1480obus[temp_w*1 +:temp_w];
assign v1480ibus[data_w*1 +:data_w] = c328obus[data_w*4 +:data_w];
assign c328ibus[temp_w*5 +:temp_w] = v1576obus[temp_w*0 +:temp_w];
assign v1576ibus[data_w*0 +:data_w] = c328obus[data_w*5 +:data_w];
assign c329ibus[temp_w*0 +:temp_w] = v6obus[temp_w*0 +:temp_w];
assign v6ibus[data_w*0 +:data_w] = c329obus[data_w*0 +:data_w];
assign c329ibus[temp_w*1 +:temp_w] = v280obus[temp_w*1 +:temp_w];
assign v280ibus[data_w*1 +:data_w] = c329obus[data_w*1 +:data_w];
assign c329ibus[temp_w*2 +:temp_w] = v778obus[temp_w*1 +:temp_w];
assign v778ibus[data_w*1 +:data_w] = c329obus[data_w*2 +:data_w];
assign c329ibus[temp_w*3 +:temp_w] = v930obus[temp_w*1 +:temp_w];
assign v930ibus[data_w*1 +:data_w] = c329obus[data_w*3 +:data_w];
assign c329ibus[temp_w*4 +:temp_w] = v1481obus[temp_w*1 +:temp_w];
assign v1481ibus[data_w*1 +:data_w] = c329obus[data_w*4 +:data_w];
assign c329ibus[temp_w*5 +:temp_w] = v1577obus[temp_w*0 +:temp_w];
assign v1577ibus[data_w*0 +:data_w] = c329obus[data_w*5 +:data_w];
assign c330ibus[temp_w*0 +:temp_w] = v7obus[temp_w*0 +:temp_w];
assign v7ibus[data_w*0 +:data_w] = c330obus[data_w*0 +:data_w];
assign c330ibus[temp_w*1 +:temp_w] = v281obus[temp_w*1 +:temp_w];
assign v281ibus[data_w*1 +:data_w] = c330obus[data_w*1 +:data_w];
assign c330ibus[temp_w*2 +:temp_w] = v779obus[temp_w*1 +:temp_w];
assign v779ibus[data_w*1 +:data_w] = c330obus[data_w*2 +:data_w];
assign c330ibus[temp_w*3 +:temp_w] = v931obus[temp_w*1 +:temp_w];
assign v931ibus[data_w*1 +:data_w] = c330obus[data_w*3 +:data_w];
assign c330ibus[temp_w*4 +:temp_w] = v1482obus[temp_w*1 +:temp_w];
assign v1482ibus[data_w*1 +:data_w] = c330obus[data_w*4 +:data_w];
assign c330ibus[temp_w*5 +:temp_w] = v1578obus[temp_w*0 +:temp_w];
assign v1578ibus[data_w*0 +:data_w] = c330obus[data_w*5 +:data_w];
assign c331ibus[temp_w*0 +:temp_w] = v8obus[temp_w*0 +:temp_w];
assign v8ibus[data_w*0 +:data_w] = c331obus[data_w*0 +:data_w];
assign c331ibus[temp_w*1 +:temp_w] = v282obus[temp_w*1 +:temp_w];
assign v282ibus[data_w*1 +:data_w] = c331obus[data_w*1 +:data_w];
assign c331ibus[temp_w*2 +:temp_w] = v780obus[temp_w*1 +:temp_w];
assign v780ibus[data_w*1 +:data_w] = c331obus[data_w*2 +:data_w];
assign c331ibus[temp_w*3 +:temp_w] = v932obus[temp_w*1 +:temp_w];
assign v932ibus[data_w*1 +:data_w] = c331obus[data_w*3 +:data_w];
assign c331ibus[temp_w*4 +:temp_w] = v1483obus[temp_w*1 +:temp_w];
assign v1483ibus[data_w*1 +:data_w] = c331obus[data_w*4 +:data_w];
assign c331ibus[temp_w*5 +:temp_w] = v1579obus[temp_w*0 +:temp_w];
assign v1579ibus[data_w*0 +:data_w] = c331obus[data_w*5 +:data_w];
assign c332ibus[temp_w*0 +:temp_w] = v9obus[temp_w*0 +:temp_w];
assign v9ibus[data_w*0 +:data_w] = c332obus[data_w*0 +:data_w];
assign c332ibus[temp_w*1 +:temp_w] = v283obus[temp_w*1 +:temp_w];
assign v283ibus[data_w*1 +:data_w] = c332obus[data_w*1 +:data_w];
assign c332ibus[temp_w*2 +:temp_w] = v781obus[temp_w*1 +:temp_w];
assign v781ibus[data_w*1 +:data_w] = c332obus[data_w*2 +:data_w];
assign c332ibus[temp_w*3 +:temp_w] = v933obus[temp_w*1 +:temp_w];
assign v933ibus[data_w*1 +:data_w] = c332obus[data_w*3 +:data_w];
assign c332ibus[temp_w*4 +:temp_w] = v1484obus[temp_w*1 +:temp_w];
assign v1484ibus[data_w*1 +:data_w] = c332obus[data_w*4 +:data_w];
assign c332ibus[temp_w*5 +:temp_w] = v1580obus[temp_w*0 +:temp_w];
assign v1580ibus[data_w*0 +:data_w] = c332obus[data_w*5 +:data_w];
assign c333ibus[temp_w*0 +:temp_w] = v10obus[temp_w*0 +:temp_w];
assign v10ibus[data_w*0 +:data_w] = c333obus[data_w*0 +:data_w];
assign c333ibus[temp_w*1 +:temp_w] = v284obus[temp_w*1 +:temp_w];
assign v284ibus[data_w*1 +:data_w] = c333obus[data_w*1 +:data_w];
assign c333ibus[temp_w*2 +:temp_w] = v782obus[temp_w*1 +:temp_w];
assign v782ibus[data_w*1 +:data_w] = c333obus[data_w*2 +:data_w];
assign c333ibus[temp_w*3 +:temp_w] = v934obus[temp_w*1 +:temp_w];
assign v934ibus[data_w*1 +:data_w] = c333obus[data_w*3 +:data_w];
assign c333ibus[temp_w*4 +:temp_w] = v1485obus[temp_w*1 +:temp_w];
assign v1485ibus[data_w*1 +:data_w] = c333obus[data_w*4 +:data_w];
assign c333ibus[temp_w*5 +:temp_w] = v1581obus[temp_w*0 +:temp_w];
assign v1581ibus[data_w*0 +:data_w] = c333obus[data_w*5 +:data_w];
assign c334ibus[temp_w*0 +:temp_w] = v11obus[temp_w*0 +:temp_w];
assign v11ibus[data_w*0 +:data_w] = c334obus[data_w*0 +:data_w];
assign c334ibus[temp_w*1 +:temp_w] = v285obus[temp_w*1 +:temp_w];
assign v285ibus[data_w*1 +:data_w] = c334obus[data_w*1 +:data_w];
assign c334ibus[temp_w*2 +:temp_w] = v783obus[temp_w*1 +:temp_w];
assign v783ibus[data_w*1 +:data_w] = c334obus[data_w*2 +:data_w];
assign c334ibus[temp_w*3 +:temp_w] = v935obus[temp_w*1 +:temp_w];
assign v935ibus[data_w*1 +:data_w] = c334obus[data_w*3 +:data_w];
assign c334ibus[temp_w*4 +:temp_w] = v1486obus[temp_w*1 +:temp_w];
assign v1486ibus[data_w*1 +:data_w] = c334obus[data_w*4 +:data_w];
assign c334ibus[temp_w*5 +:temp_w] = v1582obus[temp_w*0 +:temp_w];
assign v1582ibus[data_w*0 +:data_w] = c334obus[data_w*5 +:data_w];
assign c335ibus[temp_w*0 +:temp_w] = v12obus[temp_w*0 +:temp_w];
assign v12ibus[data_w*0 +:data_w] = c335obus[data_w*0 +:data_w];
assign c335ibus[temp_w*1 +:temp_w] = v286obus[temp_w*1 +:temp_w];
assign v286ibus[data_w*1 +:data_w] = c335obus[data_w*1 +:data_w];
assign c335ibus[temp_w*2 +:temp_w] = v784obus[temp_w*1 +:temp_w];
assign v784ibus[data_w*1 +:data_w] = c335obus[data_w*2 +:data_w];
assign c335ibus[temp_w*3 +:temp_w] = v936obus[temp_w*1 +:temp_w];
assign v936ibus[data_w*1 +:data_w] = c335obus[data_w*3 +:data_w];
assign c335ibus[temp_w*4 +:temp_w] = v1487obus[temp_w*1 +:temp_w];
assign v1487ibus[data_w*1 +:data_w] = c335obus[data_w*4 +:data_w];
assign c335ibus[temp_w*5 +:temp_w] = v1583obus[temp_w*0 +:temp_w];
assign v1583ibus[data_w*0 +:data_w] = c335obus[data_w*5 +:data_w];
assign c336ibus[temp_w*0 +:temp_w] = v13obus[temp_w*0 +:temp_w];
assign v13ibus[data_w*0 +:data_w] = c336obus[data_w*0 +:data_w];
assign c336ibus[temp_w*1 +:temp_w] = v287obus[temp_w*1 +:temp_w];
assign v287ibus[data_w*1 +:data_w] = c336obus[data_w*1 +:data_w];
assign c336ibus[temp_w*2 +:temp_w] = v785obus[temp_w*1 +:temp_w];
assign v785ibus[data_w*1 +:data_w] = c336obus[data_w*2 +:data_w];
assign c336ibus[temp_w*3 +:temp_w] = v937obus[temp_w*1 +:temp_w];
assign v937ibus[data_w*1 +:data_w] = c336obus[data_w*3 +:data_w];
assign c336ibus[temp_w*4 +:temp_w] = v1488obus[temp_w*1 +:temp_w];
assign v1488ibus[data_w*1 +:data_w] = c336obus[data_w*4 +:data_w];
assign c336ibus[temp_w*5 +:temp_w] = v1584obus[temp_w*0 +:temp_w];
assign v1584ibus[data_w*0 +:data_w] = c336obus[data_w*5 +:data_w];
assign c337ibus[temp_w*0 +:temp_w] = v14obus[temp_w*0 +:temp_w];
assign v14ibus[data_w*0 +:data_w] = c337obus[data_w*0 +:data_w];
assign c337ibus[temp_w*1 +:temp_w] = v192obus[temp_w*1 +:temp_w];
assign v192ibus[data_w*1 +:data_w] = c337obus[data_w*1 +:data_w];
assign c337ibus[temp_w*2 +:temp_w] = v786obus[temp_w*1 +:temp_w];
assign v786ibus[data_w*1 +:data_w] = c337obus[data_w*2 +:data_w];
assign c337ibus[temp_w*3 +:temp_w] = v938obus[temp_w*1 +:temp_w];
assign v938ibus[data_w*1 +:data_w] = c337obus[data_w*3 +:data_w];
assign c337ibus[temp_w*4 +:temp_w] = v1489obus[temp_w*1 +:temp_w];
assign v1489ibus[data_w*1 +:data_w] = c337obus[data_w*4 +:data_w];
assign c337ibus[temp_w*5 +:temp_w] = v1585obus[temp_w*0 +:temp_w];
assign v1585ibus[data_w*0 +:data_w] = c337obus[data_w*5 +:data_w];
assign c338ibus[temp_w*0 +:temp_w] = v15obus[temp_w*0 +:temp_w];
assign v15ibus[data_w*0 +:data_w] = c338obus[data_w*0 +:data_w];
assign c338ibus[temp_w*1 +:temp_w] = v193obus[temp_w*1 +:temp_w];
assign v193ibus[data_w*1 +:data_w] = c338obus[data_w*1 +:data_w];
assign c338ibus[temp_w*2 +:temp_w] = v787obus[temp_w*1 +:temp_w];
assign v787ibus[data_w*1 +:data_w] = c338obus[data_w*2 +:data_w];
assign c338ibus[temp_w*3 +:temp_w] = v939obus[temp_w*1 +:temp_w];
assign v939ibus[data_w*1 +:data_w] = c338obus[data_w*3 +:data_w];
assign c338ibus[temp_w*4 +:temp_w] = v1490obus[temp_w*1 +:temp_w];
assign v1490ibus[data_w*1 +:data_w] = c338obus[data_w*4 +:data_w];
assign c338ibus[temp_w*5 +:temp_w] = v1586obus[temp_w*0 +:temp_w];
assign v1586ibus[data_w*0 +:data_w] = c338obus[data_w*5 +:data_w];
assign c339ibus[temp_w*0 +:temp_w] = v16obus[temp_w*0 +:temp_w];
assign v16ibus[data_w*0 +:data_w] = c339obus[data_w*0 +:data_w];
assign c339ibus[temp_w*1 +:temp_w] = v194obus[temp_w*1 +:temp_w];
assign v194ibus[data_w*1 +:data_w] = c339obus[data_w*1 +:data_w];
assign c339ibus[temp_w*2 +:temp_w] = v788obus[temp_w*1 +:temp_w];
assign v788ibus[data_w*1 +:data_w] = c339obus[data_w*2 +:data_w];
assign c339ibus[temp_w*3 +:temp_w] = v940obus[temp_w*1 +:temp_w];
assign v940ibus[data_w*1 +:data_w] = c339obus[data_w*3 +:data_w];
assign c339ibus[temp_w*4 +:temp_w] = v1491obus[temp_w*1 +:temp_w];
assign v1491ibus[data_w*1 +:data_w] = c339obus[data_w*4 +:data_w];
assign c339ibus[temp_w*5 +:temp_w] = v1587obus[temp_w*0 +:temp_w];
assign v1587ibus[data_w*0 +:data_w] = c339obus[data_w*5 +:data_w];
assign c340ibus[temp_w*0 +:temp_w] = v17obus[temp_w*0 +:temp_w];
assign v17ibus[data_w*0 +:data_w] = c340obus[data_w*0 +:data_w];
assign c340ibus[temp_w*1 +:temp_w] = v195obus[temp_w*1 +:temp_w];
assign v195ibus[data_w*1 +:data_w] = c340obus[data_w*1 +:data_w];
assign c340ibus[temp_w*2 +:temp_w] = v789obus[temp_w*1 +:temp_w];
assign v789ibus[data_w*1 +:data_w] = c340obus[data_w*2 +:data_w];
assign c340ibus[temp_w*3 +:temp_w] = v941obus[temp_w*1 +:temp_w];
assign v941ibus[data_w*1 +:data_w] = c340obus[data_w*3 +:data_w];
assign c340ibus[temp_w*4 +:temp_w] = v1492obus[temp_w*1 +:temp_w];
assign v1492ibus[data_w*1 +:data_w] = c340obus[data_w*4 +:data_w];
assign c340ibus[temp_w*5 +:temp_w] = v1588obus[temp_w*0 +:temp_w];
assign v1588ibus[data_w*0 +:data_w] = c340obus[data_w*5 +:data_w];
assign c341ibus[temp_w*0 +:temp_w] = v18obus[temp_w*0 +:temp_w];
assign v18ibus[data_w*0 +:data_w] = c341obus[data_w*0 +:data_w];
assign c341ibus[temp_w*1 +:temp_w] = v196obus[temp_w*1 +:temp_w];
assign v196ibus[data_w*1 +:data_w] = c341obus[data_w*1 +:data_w];
assign c341ibus[temp_w*2 +:temp_w] = v790obus[temp_w*1 +:temp_w];
assign v790ibus[data_w*1 +:data_w] = c341obus[data_w*2 +:data_w];
assign c341ibus[temp_w*3 +:temp_w] = v942obus[temp_w*1 +:temp_w];
assign v942ibus[data_w*1 +:data_w] = c341obus[data_w*3 +:data_w];
assign c341ibus[temp_w*4 +:temp_w] = v1493obus[temp_w*1 +:temp_w];
assign v1493ibus[data_w*1 +:data_w] = c341obus[data_w*4 +:data_w];
assign c341ibus[temp_w*5 +:temp_w] = v1589obus[temp_w*0 +:temp_w];
assign v1589ibus[data_w*0 +:data_w] = c341obus[data_w*5 +:data_w];
assign c342ibus[temp_w*0 +:temp_w] = v19obus[temp_w*0 +:temp_w];
assign v19ibus[data_w*0 +:data_w] = c342obus[data_w*0 +:data_w];
assign c342ibus[temp_w*1 +:temp_w] = v197obus[temp_w*1 +:temp_w];
assign v197ibus[data_w*1 +:data_w] = c342obus[data_w*1 +:data_w];
assign c342ibus[temp_w*2 +:temp_w] = v791obus[temp_w*1 +:temp_w];
assign v791ibus[data_w*1 +:data_w] = c342obus[data_w*2 +:data_w];
assign c342ibus[temp_w*3 +:temp_w] = v943obus[temp_w*1 +:temp_w];
assign v943ibus[data_w*1 +:data_w] = c342obus[data_w*3 +:data_w];
assign c342ibus[temp_w*4 +:temp_w] = v1494obus[temp_w*1 +:temp_w];
assign v1494ibus[data_w*1 +:data_w] = c342obus[data_w*4 +:data_w];
assign c342ibus[temp_w*5 +:temp_w] = v1590obus[temp_w*0 +:temp_w];
assign v1590ibus[data_w*0 +:data_w] = c342obus[data_w*5 +:data_w];
assign c343ibus[temp_w*0 +:temp_w] = v20obus[temp_w*0 +:temp_w];
assign v20ibus[data_w*0 +:data_w] = c343obus[data_w*0 +:data_w];
assign c343ibus[temp_w*1 +:temp_w] = v198obus[temp_w*1 +:temp_w];
assign v198ibus[data_w*1 +:data_w] = c343obus[data_w*1 +:data_w];
assign c343ibus[temp_w*2 +:temp_w] = v792obus[temp_w*1 +:temp_w];
assign v792ibus[data_w*1 +:data_w] = c343obus[data_w*2 +:data_w];
assign c343ibus[temp_w*3 +:temp_w] = v944obus[temp_w*1 +:temp_w];
assign v944ibus[data_w*1 +:data_w] = c343obus[data_w*3 +:data_w];
assign c343ibus[temp_w*4 +:temp_w] = v1495obus[temp_w*1 +:temp_w];
assign v1495ibus[data_w*1 +:data_w] = c343obus[data_w*4 +:data_w];
assign c343ibus[temp_w*5 +:temp_w] = v1591obus[temp_w*0 +:temp_w];
assign v1591ibus[data_w*0 +:data_w] = c343obus[data_w*5 +:data_w];
assign c344ibus[temp_w*0 +:temp_w] = v21obus[temp_w*0 +:temp_w];
assign v21ibus[data_w*0 +:data_w] = c344obus[data_w*0 +:data_w];
assign c344ibus[temp_w*1 +:temp_w] = v199obus[temp_w*1 +:temp_w];
assign v199ibus[data_w*1 +:data_w] = c344obus[data_w*1 +:data_w];
assign c344ibus[temp_w*2 +:temp_w] = v793obus[temp_w*1 +:temp_w];
assign v793ibus[data_w*1 +:data_w] = c344obus[data_w*2 +:data_w];
assign c344ibus[temp_w*3 +:temp_w] = v945obus[temp_w*1 +:temp_w];
assign v945ibus[data_w*1 +:data_w] = c344obus[data_w*3 +:data_w];
assign c344ibus[temp_w*4 +:temp_w] = v1496obus[temp_w*1 +:temp_w];
assign v1496ibus[data_w*1 +:data_w] = c344obus[data_w*4 +:data_w];
assign c344ibus[temp_w*5 +:temp_w] = v1592obus[temp_w*0 +:temp_w];
assign v1592ibus[data_w*0 +:data_w] = c344obus[data_w*5 +:data_w];
assign c345ibus[temp_w*0 +:temp_w] = v22obus[temp_w*0 +:temp_w];
assign v22ibus[data_w*0 +:data_w] = c345obus[data_w*0 +:data_w];
assign c345ibus[temp_w*1 +:temp_w] = v200obus[temp_w*1 +:temp_w];
assign v200ibus[data_w*1 +:data_w] = c345obus[data_w*1 +:data_w];
assign c345ibus[temp_w*2 +:temp_w] = v794obus[temp_w*1 +:temp_w];
assign v794ibus[data_w*1 +:data_w] = c345obus[data_w*2 +:data_w];
assign c345ibus[temp_w*3 +:temp_w] = v946obus[temp_w*1 +:temp_w];
assign v946ibus[data_w*1 +:data_w] = c345obus[data_w*3 +:data_w];
assign c345ibus[temp_w*4 +:temp_w] = v1497obus[temp_w*1 +:temp_w];
assign v1497ibus[data_w*1 +:data_w] = c345obus[data_w*4 +:data_w];
assign c345ibus[temp_w*5 +:temp_w] = v1593obus[temp_w*0 +:temp_w];
assign v1593ibus[data_w*0 +:data_w] = c345obus[data_w*5 +:data_w];
assign c346ibus[temp_w*0 +:temp_w] = v23obus[temp_w*0 +:temp_w];
assign v23ibus[data_w*0 +:data_w] = c346obus[data_w*0 +:data_w];
assign c346ibus[temp_w*1 +:temp_w] = v201obus[temp_w*1 +:temp_w];
assign v201ibus[data_w*1 +:data_w] = c346obus[data_w*1 +:data_w];
assign c346ibus[temp_w*2 +:temp_w] = v795obus[temp_w*1 +:temp_w];
assign v795ibus[data_w*1 +:data_w] = c346obus[data_w*2 +:data_w];
assign c346ibus[temp_w*3 +:temp_w] = v947obus[temp_w*1 +:temp_w];
assign v947ibus[data_w*1 +:data_w] = c346obus[data_w*3 +:data_w];
assign c346ibus[temp_w*4 +:temp_w] = v1498obus[temp_w*1 +:temp_w];
assign v1498ibus[data_w*1 +:data_w] = c346obus[data_w*4 +:data_w];
assign c346ibus[temp_w*5 +:temp_w] = v1594obus[temp_w*0 +:temp_w];
assign v1594ibus[data_w*0 +:data_w] = c346obus[data_w*5 +:data_w];
assign c347ibus[temp_w*0 +:temp_w] = v24obus[temp_w*0 +:temp_w];
assign v24ibus[data_w*0 +:data_w] = c347obus[data_w*0 +:data_w];
assign c347ibus[temp_w*1 +:temp_w] = v202obus[temp_w*1 +:temp_w];
assign v202ibus[data_w*1 +:data_w] = c347obus[data_w*1 +:data_w];
assign c347ibus[temp_w*2 +:temp_w] = v796obus[temp_w*1 +:temp_w];
assign v796ibus[data_w*1 +:data_w] = c347obus[data_w*2 +:data_w];
assign c347ibus[temp_w*3 +:temp_w] = v948obus[temp_w*1 +:temp_w];
assign v948ibus[data_w*1 +:data_w] = c347obus[data_w*3 +:data_w];
assign c347ibus[temp_w*4 +:temp_w] = v1499obus[temp_w*1 +:temp_w];
assign v1499ibus[data_w*1 +:data_w] = c347obus[data_w*4 +:data_w];
assign c347ibus[temp_w*5 +:temp_w] = v1595obus[temp_w*0 +:temp_w];
assign v1595ibus[data_w*0 +:data_w] = c347obus[data_w*5 +:data_w];
assign c348ibus[temp_w*0 +:temp_w] = v25obus[temp_w*0 +:temp_w];
assign v25ibus[data_w*0 +:data_w] = c348obus[data_w*0 +:data_w];
assign c348ibus[temp_w*1 +:temp_w] = v203obus[temp_w*1 +:temp_w];
assign v203ibus[data_w*1 +:data_w] = c348obus[data_w*1 +:data_w];
assign c348ibus[temp_w*2 +:temp_w] = v797obus[temp_w*1 +:temp_w];
assign v797ibus[data_w*1 +:data_w] = c348obus[data_w*2 +:data_w];
assign c348ibus[temp_w*3 +:temp_w] = v949obus[temp_w*1 +:temp_w];
assign v949ibus[data_w*1 +:data_w] = c348obus[data_w*3 +:data_w];
assign c348ibus[temp_w*4 +:temp_w] = v1500obus[temp_w*1 +:temp_w];
assign v1500ibus[data_w*1 +:data_w] = c348obus[data_w*4 +:data_w];
assign c348ibus[temp_w*5 +:temp_w] = v1596obus[temp_w*0 +:temp_w];
assign v1596ibus[data_w*0 +:data_w] = c348obus[data_w*5 +:data_w];
assign c349ibus[temp_w*0 +:temp_w] = v26obus[temp_w*0 +:temp_w];
assign v26ibus[data_w*0 +:data_w] = c349obus[data_w*0 +:data_w];
assign c349ibus[temp_w*1 +:temp_w] = v204obus[temp_w*1 +:temp_w];
assign v204ibus[data_w*1 +:data_w] = c349obus[data_w*1 +:data_w];
assign c349ibus[temp_w*2 +:temp_w] = v798obus[temp_w*1 +:temp_w];
assign v798ibus[data_w*1 +:data_w] = c349obus[data_w*2 +:data_w];
assign c349ibus[temp_w*3 +:temp_w] = v950obus[temp_w*1 +:temp_w];
assign v950ibus[data_w*1 +:data_w] = c349obus[data_w*3 +:data_w];
assign c349ibus[temp_w*4 +:temp_w] = v1501obus[temp_w*1 +:temp_w];
assign v1501ibus[data_w*1 +:data_w] = c349obus[data_w*4 +:data_w];
assign c349ibus[temp_w*5 +:temp_w] = v1597obus[temp_w*0 +:temp_w];
assign v1597ibus[data_w*0 +:data_w] = c349obus[data_w*5 +:data_w];
assign c350ibus[temp_w*0 +:temp_w] = v27obus[temp_w*0 +:temp_w];
assign v27ibus[data_w*0 +:data_w] = c350obus[data_w*0 +:data_w];
assign c350ibus[temp_w*1 +:temp_w] = v205obus[temp_w*1 +:temp_w];
assign v205ibus[data_w*1 +:data_w] = c350obus[data_w*1 +:data_w];
assign c350ibus[temp_w*2 +:temp_w] = v799obus[temp_w*1 +:temp_w];
assign v799ibus[data_w*1 +:data_w] = c350obus[data_w*2 +:data_w];
assign c350ibus[temp_w*3 +:temp_w] = v951obus[temp_w*1 +:temp_w];
assign v951ibus[data_w*1 +:data_w] = c350obus[data_w*3 +:data_w];
assign c350ibus[temp_w*4 +:temp_w] = v1502obus[temp_w*1 +:temp_w];
assign v1502ibus[data_w*1 +:data_w] = c350obus[data_w*4 +:data_w];
assign c350ibus[temp_w*5 +:temp_w] = v1598obus[temp_w*0 +:temp_w];
assign v1598ibus[data_w*0 +:data_w] = c350obus[data_w*5 +:data_w];
assign c351ibus[temp_w*0 +:temp_w] = v28obus[temp_w*0 +:temp_w];
assign v28ibus[data_w*0 +:data_w] = c351obus[data_w*0 +:data_w];
assign c351ibus[temp_w*1 +:temp_w] = v206obus[temp_w*1 +:temp_w];
assign v206ibus[data_w*1 +:data_w] = c351obus[data_w*1 +:data_w];
assign c351ibus[temp_w*2 +:temp_w] = v800obus[temp_w*1 +:temp_w];
assign v800ibus[data_w*1 +:data_w] = c351obus[data_w*2 +:data_w];
assign c351ibus[temp_w*3 +:temp_w] = v952obus[temp_w*1 +:temp_w];
assign v952ibus[data_w*1 +:data_w] = c351obus[data_w*3 +:data_w];
assign c351ibus[temp_w*4 +:temp_w] = v1503obus[temp_w*1 +:temp_w];
assign v1503ibus[data_w*1 +:data_w] = c351obus[data_w*4 +:data_w];
assign c351ibus[temp_w*5 +:temp_w] = v1599obus[temp_w*0 +:temp_w];
assign v1599ibus[data_w*0 +:data_w] = c351obus[data_w*5 +:data_w];
assign c352ibus[temp_w*0 +:temp_w] = v29obus[temp_w*0 +:temp_w];
assign v29ibus[data_w*0 +:data_w] = c352obus[data_w*0 +:data_w];
assign c352ibus[temp_w*1 +:temp_w] = v207obus[temp_w*1 +:temp_w];
assign v207ibus[data_w*1 +:data_w] = c352obus[data_w*1 +:data_w];
assign c352ibus[temp_w*2 +:temp_w] = v801obus[temp_w*1 +:temp_w];
assign v801ibus[data_w*1 +:data_w] = c352obus[data_w*2 +:data_w];
assign c352ibus[temp_w*3 +:temp_w] = v953obus[temp_w*1 +:temp_w];
assign v953ibus[data_w*1 +:data_w] = c352obus[data_w*3 +:data_w];
assign c352ibus[temp_w*4 +:temp_w] = v1504obus[temp_w*1 +:temp_w];
assign v1504ibus[data_w*1 +:data_w] = c352obus[data_w*4 +:data_w];
assign c352ibus[temp_w*5 +:temp_w] = v1600obus[temp_w*0 +:temp_w];
assign v1600ibus[data_w*0 +:data_w] = c352obus[data_w*5 +:data_w];
assign c353ibus[temp_w*0 +:temp_w] = v30obus[temp_w*0 +:temp_w];
assign v30ibus[data_w*0 +:data_w] = c353obus[data_w*0 +:data_w];
assign c353ibus[temp_w*1 +:temp_w] = v208obus[temp_w*1 +:temp_w];
assign v208ibus[data_w*1 +:data_w] = c353obus[data_w*1 +:data_w];
assign c353ibus[temp_w*2 +:temp_w] = v802obus[temp_w*1 +:temp_w];
assign v802ibus[data_w*1 +:data_w] = c353obus[data_w*2 +:data_w];
assign c353ibus[temp_w*3 +:temp_w] = v954obus[temp_w*1 +:temp_w];
assign v954ibus[data_w*1 +:data_w] = c353obus[data_w*3 +:data_w];
assign c353ibus[temp_w*4 +:temp_w] = v1505obus[temp_w*1 +:temp_w];
assign v1505ibus[data_w*1 +:data_w] = c353obus[data_w*4 +:data_w];
assign c353ibus[temp_w*5 +:temp_w] = v1601obus[temp_w*0 +:temp_w];
assign v1601ibus[data_w*0 +:data_w] = c353obus[data_w*5 +:data_w];
assign c354ibus[temp_w*0 +:temp_w] = v31obus[temp_w*0 +:temp_w];
assign v31ibus[data_w*0 +:data_w] = c354obus[data_w*0 +:data_w];
assign c354ibus[temp_w*1 +:temp_w] = v209obus[temp_w*1 +:temp_w];
assign v209ibus[data_w*1 +:data_w] = c354obus[data_w*1 +:data_w];
assign c354ibus[temp_w*2 +:temp_w] = v803obus[temp_w*1 +:temp_w];
assign v803ibus[data_w*1 +:data_w] = c354obus[data_w*2 +:data_w];
assign c354ibus[temp_w*3 +:temp_w] = v955obus[temp_w*1 +:temp_w];
assign v955ibus[data_w*1 +:data_w] = c354obus[data_w*3 +:data_w];
assign c354ibus[temp_w*4 +:temp_w] = v1506obus[temp_w*1 +:temp_w];
assign v1506ibus[data_w*1 +:data_w] = c354obus[data_w*4 +:data_w];
assign c354ibus[temp_w*5 +:temp_w] = v1602obus[temp_w*0 +:temp_w];
assign v1602ibus[data_w*0 +:data_w] = c354obus[data_w*5 +:data_w];
assign c355ibus[temp_w*0 +:temp_w] = v32obus[temp_w*0 +:temp_w];
assign v32ibus[data_w*0 +:data_w] = c355obus[data_w*0 +:data_w];
assign c355ibus[temp_w*1 +:temp_w] = v210obus[temp_w*1 +:temp_w];
assign v210ibus[data_w*1 +:data_w] = c355obus[data_w*1 +:data_w];
assign c355ibus[temp_w*2 +:temp_w] = v804obus[temp_w*1 +:temp_w];
assign v804ibus[data_w*1 +:data_w] = c355obus[data_w*2 +:data_w];
assign c355ibus[temp_w*3 +:temp_w] = v956obus[temp_w*1 +:temp_w];
assign v956ibus[data_w*1 +:data_w] = c355obus[data_w*3 +:data_w];
assign c355ibus[temp_w*4 +:temp_w] = v1507obus[temp_w*1 +:temp_w];
assign v1507ibus[data_w*1 +:data_w] = c355obus[data_w*4 +:data_w];
assign c355ibus[temp_w*5 +:temp_w] = v1603obus[temp_w*0 +:temp_w];
assign v1603ibus[data_w*0 +:data_w] = c355obus[data_w*5 +:data_w];
assign c356ibus[temp_w*0 +:temp_w] = v33obus[temp_w*0 +:temp_w];
assign v33ibus[data_w*0 +:data_w] = c356obus[data_w*0 +:data_w];
assign c356ibus[temp_w*1 +:temp_w] = v211obus[temp_w*1 +:temp_w];
assign v211ibus[data_w*1 +:data_w] = c356obus[data_w*1 +:data_w];
assign c356ibus[temp_w*2 +:temp_w] = v805obus[temp_w*1 +:temp_w];
assign v805ibus[data_w*1 +:data_w] = c356obus[data_w*2 +:data_w];
assign c356ibus[temp_w*3 +:temp_w] = v957obus[temp_w*1 +:temp_w];
assign v957ibus[data_w*1 +:data_w] = c356obus[data_w*3 +:data_w];
assign c356ibus[temp_w*4 +:temp_w] = v1508obus[temp_w*1 +:temp_w];
assign v1508ibus[data_w*1 +:data_w] = c356obus[data_w*4 +:data_w];
assign c356ibus[temp_w*5 +:temp_w] = v1604obus[temp_w*0 +:temp_w];
assign v1604ibus[data_w*0 +:data_w] = c356obus[data_w*5 +:data_w];
assign c357ibus[temp_w*0 +:temp_w] = v34obus[temp_w*0 +:temp_w];
assign v34ibus[data_w*0 +:data_w] = c357obus[data_w*0 +:data_w];
assign c357ibus[temp_w*1 +:temp_w] = v212obus[temp_w*1 +:temp_w];
assign v212ibus[data_w*1 +:data_w] = c357obus[data_w*1 +:data_w];
assign c357ibus[temp_w*2 +:temp_w] = v806obus[temp_w*1 +:temp_w];
assign v806ibus[data_w*1 +:data_w] = c357obus[data_w*2 +:data_w];
assign c357ibus[temp_w*3 +:temp_w] = v958obus[temp_w*1 +:temp_w];
assign v958ibus[data_w*1 +:data_w] = c357obus[data_w*3 +:data_w];
assign c357ibus[temp_w*4 +:temp_w] = v1509obus[temp_w*1 +:temp_w];
assign v1509ibus[data_w*1 +:data_w] = c357obus[data_w*4 +:data_w];
assign c357ibus[temp_w*5 +:temp_w] = v1605obus[temp_w*0 +:temp_w];
assign v1605ibus[data_w*0 +:data_w] = c357obus[data_w*5 +:data_w];
assign c358ibus[temp_w*0 +:temp_w] = v35obus[temp_w*0 +:temp_w];
assign v35ibus[data_w*0 +:data_w] = c358obus[data_w*0 +:data_w];
assign c358ibus[temp_w*1 +:temp_w] = v213obus[temp_w*1 +:temp_w];
assign v213ibus[data_w*1 +:data_w] = c358obus[data_w*1 +:data_w];
assign c358ibus[temp_w*2 +:temp_w] = v807obus[temp_w*1 +:temp_w];
assign v807ibus[data_w*1 +:data_w] = c358obus[data_w*2 +:data_w];
assign c358ibus[temp_w*3 +:temp_w] = v959obus[temp_w*1 +:temp_w];
assign v959ibus[data_w*1 +:data_w] = c358obus[data_w*3 +:data_w];
assign c358ibus[temp_w*4 +:temp_w] = v1510obus[temp_w*1 +:temp_w];
assign v1510ibus[data_w*1 +:data_w] = c358obus[data_w*4 +:data_w];
assign c358ibus[temp_w*5 +:temp_w] = v1606obus[temp_w*0 +:temp_w];
assign v1606ibus[data_w*0 +:data_w] = c358obus[data_w*5 +:data_w];
assign c359ibus[temp_w*0 +:temp_w] = v36obus[temp_w*0 +:temp_w];
assign v36ibus[data_w*0 +:data_w] = c359obus[data_w*0 +:data_w];
assign c359ibus[temp_w*1 +:temp_w] = v214obus[temp_w*1 +:temp_w];
assign v214ibus[data_w*1 +:data_w] = c359obus[data_w*1 +:data_w];
assign c359ibus[temp_w*2 +:temp_w] = v808obus[temp_w*1 +:temp_w];
assign v808ibus[data_w*1 +:data_w] = c359obus[data_w*2 +:data_w];
assign c359ibus[temp_w*3 +:temp_w] = v864obus[temp_w*1 +:temp_w];
assign v864ibus[data_w*1 +:data_w] = c359obus[data_w*3 +:data_w];
assign c359ibus[temp_w*4 +:temp_w] = v1511obus[temp_w*1 +:temp_w];
assign v1511ibus[data_w*1 +:data_w] = c359obus[data_w*4 +:data_w];
assign c359ibus[temp_w*5 +:temp_w] = v1607obus[temp_w*0 +:temp_w];
assign v1607ibus[data_w*0 +:data_w] = c359obus[data_w*5 +:data_w];
assign c360ibus[temp_w*0 +:temp_w] = v37obus[temp_w*0 +:temp_w];
assign v37ibus[data_w*0 +:data_w] = c360obus[data_w*0 +:data_w];
assign c360ibus[temp_w*1 +:temp_w] = v215obus[temp_w*1 +:temp_w];
assign v215ibus[data_w*1 +:data_w] = c360obus[data_w*1 +:data_w];
assign c360ibus[temp_w*2 +:temp_w] = v809obus[temp_w*1 +:temp_w];
assign v809ibus[data_w*1 +:data_w] = c360obus[data_w*2 +:data_w];
assign c360ibus[temp_w*3 +:temp_w] = v865obus[temp_w*1 +:temp_w];
assign v865ibus[data_w*1 +:data_w] = c360obus[data_w*3 +:data_w];
assign c360ibus[temp_w*4 +:temp_w] = v1512obus[temp_w*1 +:temp_w];
assign v1512ibus[data_w*1 +:data_w] = c360obus[data_w*4 +:data_w];
assign c360ibus[temp_w*5 +:temp_w] = v1608obus[temp_w*0 +:temp_w];
assign v1608ibus[data_w*0 +:data_w] = c360obus[data_w*5 +:data_w];
assign c361ibus[temp_w*0 +:temp_w] = v38obus[temp_w*0 +:temp_w];
assign v38ibus[data_w*0 +:data_w] = c361obus[data_w*0 +:data_w];
assign c361ibus[temp_w*1 +:temp_w] = v216obus[temp_w*1 +:temp_w];
assign v216ibus[data_w*1 +:data_w] = c361obus[data_w*1 +:data_w];
assign c361ibus[temp_w*2 +:temp_w] = v810obus[temp_w*1 +:temp_w];
assign v810ibus[data_w*1 +:data_w] = c361obus[data_w*2 +:data_w];
assign c361ibus[temp_w*3 +:temp_w] = v866obus[temp_w*1 +:temp_w];
assign v866ibus[data_w*1 +:data_w] = c361obus[data_w*3 +:data_w];
assign c361ibus[temp_w*4 +:temp_w] = v1513obus[temp_w*1 +:temp_w];
assign v1513ibus[data_w*1 +:data_w] = c361obus[data_w*4 +:data_w];
assign c361ibus[temp_w*5 +:temp_w] = v1609obus[temp_w*0 +:temp_w];
assign v1609ibus[data_w*0 +:data_w] = c361obus[data_w*5 +:data_w];
assign c362ibus[temp_w*0 +:temp_w] = v39obus[temp_w*0 +:temp_w];
assign v39ibus[data_w*0 +:data_w] = c362obus[data_w*0 +:data_w];
assign c362ibus[temp_w*1 +:temp_w] = v217obus[temp_w*1 +:temp_w];
assign v217ibus[data_w*1 +:data_w] = c362obus[data_w*1 +:data_w];
assign c362ibus[temp_w*2 +:temp_w] = v811obus[temp_w*1 +:temp_w];
assign v811ibus[data_w*1 +:data_w] = c362obus[data_w*2 +:data_w];
assign c362ibus[temp_w*3 +:temp_w] = v867obus[temp_w*1 +:temp_w];
assign v867ibus[data_w*1 +:data_w] = c362obus[data_w*3 +:data_w];
assign c362ibus[temp_w*4 +:temp_w] = v1514obus[temp_w*1 +:temp_w];
assign v1514ibus[data_w*1 +:data_w] = c362obus[data_w*4 +:data_w];
assign c362ibus[temp_w*5 +:temp_w] = v1610obus[temp_w*0 +:temp_w];
assign v1610ibus[data_w*0 +:data_w] = c362obus[data_w*5 +:data_w];
assign c363ibus[temp_w*0 +:temp_w] = v40obus[temp_w*0 +:temp_w];
assign v40ibus[data_w*0 +:data_w] = c363obus[data_w*0 +:data_w];
assign c363ibus[temp_w*1 +:temp_w] = v218obus[temp_w*1 +:temp_w];
assign v218ibus[data_w*1 +:data_w] = c363obus[data_w*1 +:data_w];
assign c363ibus[temp_w*2 +:temp_w] = v812obus[temp_w*1 +:temp_w];
assign v812ibus[data_w*1 +:data_w] = c363obus[data_w*2 +:data_w];
assign c363ibus[temp_w*3 +:temp_w] = v868obus[temp_w*1 +:temp_w];
assign v868ibus[data_w*1 +:data_w] = c363obus[data_w*3 +:data_w];
assign c363ibus[temp_w*4 +:temp_w] = v1515obus[temp_w*1 +:temp_w];
assign v1515ibus[data_w*1 +:data_w] = c363obus[data_w*4 +:data_w];
assign c363ibus[temp_w*5 +:temp_w] = v1611obus[temp_w*0 +:temp_w];
assign v1611ibus[data_w*0 +:data_w] = c363obus[data_w*5 +:data_w];
assign c364ibus[temp_w*0 +:temp_w] = v41obus[temp_w*0 +:temp_w];
assign v41ibus[data_w*0 +:data_w] = c364obus[data_w*0 +:data_w];
assign c364ibus[temp_w*1 +:temp_w] = v219obus[temp_w*1 +:temp_w];
assign v219ibus[data_w*1 +:data_w] = c364obus[data_w*1 +:data_w];
assign c364ibus[temp_w*2 +:temp_w] = v813obus[temp_w*1 +:temp_w];
assign v813ibus[data_w*1 +:data_w] = c364obus[data_w*2 +:data_w];
assign c364ibus[temp_w*3 +:temp_w] = v869obus[temp_w*1 +:temp_w];
assign v869ibus[data_w*1 +:data_w] = c364obus[data_w*3 +:data_w];
assign c364ibus[temp_w*4 +:temp_w] = v1516obus[temp_w*1 +:temp_w];
assign v1516ibus[data_w*1 +:data_w] = c364obus[data_w*4 +:data_w];
assign c364ibus[temp_w*5 +:temp_w] = v1612obus[temp_w*0 +:temp_w];
assign v1612ibus[data_w*0 +:data_w] = c364obus[data_w*5 +:data_w];
assign c365ibus[temp_w*0 +:temp_w] = v42obus[temp_w*0 +:temp_w];
assign v42ibus[data_w*0 +:data_w] = c365obus[data_w*0 +:data_w];
assign c365ibus[temp_w*1 +:temp_w] = v220obus[temp_w*1 +:temp_w];
assign v220ibus[data_w*1 +:data_w] = c365obus[data_w*1 +:data_w];
assign c365ibus[temp_w*2 +:temp_w] = v814obus[temp_w*1 +:temp_w];
assign v814ibus[data_w*1 +:data_w] = c365obus[data_w*2 +:data_w];
assign c365ibus[temp_w*3 +:temp_w] = v870obus[temp_w*1 +:temp_w];
assign v870ibus[data_w*1 +:data_w] = c365obus[data_w*3 +:data_w];
assign c365ibus[temp_w*4 +:temp_w] = v1517obus[temp_w*1 +:temp_w];
assign v1517ibus[data_w*1 +:data_w] = c365obus[data_w*4 +:data_w];
assign c365ibus[temp_w*5 +:temp_w] = v1613obus[temp_w*0 +:temp_w];
assign v1613ibus[data_w*0 +:data_w] = c365obus[data_w*5 +:data_w];
assign c366ibus[temp_w*0 +:temp_w] = v43obus[temp_w*0 +:temp_w];
assign v43ibus[data_w*0 +:data_w] = c366obus[data_w*0 +:data_w];
assign c366ibus[temp_w*1 +:temp_w] = v221obus[temp_w*1 +:temp_w];
assign v221ibus[data_w*1 +:data_w] = c366obus[data_w*1 +:data_w];
assign c366ibus[temp_w*2 +:temp_w] = v815obus[temp_w*1 +:temp_w];
assign v815ibus[data_w*1 +:data_w] = c366obus[data_w*2 +:data_w];
assign c366ibus[temp_w*3 +:temp_w] = v871obus[temp_w*1 +:temp_w];
assign v871ibus[data_w*1 +:data_w] = c366obus[data_w*3 +:data_w];
assign c366ibus[temp_w*4 +:temp_w] = v1518obus[temp_w*1 +:temp_w];
assign v1518ibus[data_w*1 +:data_w] = c366obus[data_w*4 +:data_w];
assign c366ibus[temp_w*5 +:temp_w] = v1614obus[temp_w*0 +:temp_w];
assign v1614ibus[data_w*0 +:data_w] = c366obus[data_w*5 +:data_w];
assign c367ibus[temp_w*0 +:temp_w] = v44obus[temp_w*0 +:temp_w];
assign v44ibus[data_w*0 +:data_w] = c367obus[data_w*0 +:data_w];
assign c367ibus[temp_w*1 +:temp_w] = v222obus[temp_w*1 +:temp_w];
assign v222ibus[data_w*1 +:data_w] = c367obus[data_w*1 +:data_w];
assign c367ibus[temp_w*2 +:temp_w] = v816obus[temp_w*1 +:temp_w];
assign v816ibus[data_w*1 +:data_w] = c367obus[data_w*2 +:data_w];
assign c367ibus[temp_w*3 +:temp_w] = v872obus[temp_w*1 +:temp_w];
assign v872ibus[data_w*1 +:data_w] = c367obus[data_w*3 +:data_w];
assign c367ibus[temp_w*4 +:temp_w] = v1519obus[temp_w*1 +:temp_w];
assign v1519ibus[data_w*1 +:data_w] = c367obus[data_w*4 +:data_w];
assign c367ibus[temp_w*5 +:temp_w] = v1615obus[temp_w*0 +:temp_w];
assign v1615ibus[data_w*0 +:data_w] = c367obus[data_w*5 +:data_w];
assign c368ibus[temp_w*0 +:temp_w] = v45obus[temp_w*0 +:temp_w];
assign v45ibus[data_w*0 +:data_w] = c368obus[data_w*0 +:data_w];
assign c368ibus[temp_w*1 +:temp_w] = v223obus[temp_w*1 +:temp_w];
assign v223ibus[data_w*1 +:data_w] = c368obus[data_w*1 +:data_w];
assign c368ibus[temp_w*2 +:temp_w] = v817obus[temp_w*1 +:temp_w];
assign v817ibus[data_w*1 +:data_w] = c368obus[data_w*2 +:data_w];
assign c368ibus[temp_w*3 +:temp_w] = v873obus[temp_w*1 +:temp_w];
assign v873ibus[data_w*1 +:data_w] = c368obus[data_w*3 +:data_w];
assign c368ibus[temp_w*4 +:temp_w] = v1520obus[temp_w*1 +:temp_w];
assign v1520ibus[data_w*1 +:data_w] = c368obus[data_w*4 +:data_w];
assign c368ibus[temp_w*5 +:temp_w] = v1616obus[temp_w*0 +:temp_w];
assign v1616ibus[data_w*0 +:data_w] = c368obus[data_w*5 +:data_w];
assign c369ibus[temp_w*0 +:temp_w] = v46obus[temp_w*0 +:temp_w];
assign v46ibus[data_w*0 +:data_w] = c369obus[data_w*0 +:data_w];
assign c369ibus[temp_w*1 +:temp_w] = v224obus[temp_w*1 +:temp_w];
assign v224ibus[data_w*1 +:data_w] = c369obus[data_w*1 +:data_w];
assign c369ibus[temp_w*2 +:temp_w] = v818obus[temp_w*1 +:temp_w];
assign v818ibus[data_w*1 +:data_w] = c369obus[data_w*2 +:data_w];
assign c369ibus[temp_w*3 +:temp_w] = v874obus[temp_w*1 +:temp_w];
assign v874ibus[data_w*1 +:data_w] = c369obus[data_w*3 +:data_w];
assign c369ibus[temp_w*4 +:temp_w] = v1521obus[temp_w*1 +:temp_w];
assign v1521ibus[data_w*1 +:data_w] = c369obus[data_w*4 +:data_w];
assign c369ibus[temp_w*5 +:temp_w] = v1617obus[temp_w*0 +:temp_w];
assign v1617ibus[data_w*0 +:data_w] = c369obus[data_w*5 +:data_w];
assign c370ibus[temp_w*0 +:temp_w] = v47obus[temp_w*0 +:temp_w];
assign v47ibus[data_w*0 +:data_w] = c370obus[data_w*0 +:data_w];
assign c370ibus[temp_w*1 +:temp_w] = v225obus[temp_w*1 +:temp_w];
assign v225ibus[data_w*1 +:data_w] = c370obus[data_w*1 +:data_w];
assign c370ibus[temp_w*2 +:temp_w] = v819obus[temp_w*1 +:temp_w];
assign v819ibus[data_w*1 +:data_w] = c370obus[data_w*2 +:data_w];
assign c370ibus[temp_w*3 +:temp_w] = v875obus[temp_w*1 +:temp_w];
assign v875ibus[data_w*1 +:data_w] = c370obus[data_w*3 +:data_w];
assign c370ibus[temp_w*4 +:temp_w] = v1522obus[temp_w*1 +:temp_w];
assign v1522ibus[data_w*1 +:data_w] = c370obus[data_w*4 +:data_w];
assign c370ibus[temp_w*5 +:temp_w] = v1618obus[temp_w*0 +:temp_w];
assign v1618ibus[data_w*0 +:data_w] = c370obus[data_w*5 +:data_w];
assign c371ibus[temp_w*0 +:temp_w] = v48obus[temp_w*0 +:temp_w];
assign v48ibus[data_w*0 +:data_w] = c371obus[data_w*0 +:data_w];
assign c371ibus[temp_w*1 +:temp_w] = v226obus[temp_w*1 +:temp_w];
assign v226ibus[data_w*1 +:data_w] = c371obus[data_w*1 +:data_w];
assign c371ibus[temp_w*2 +:temp_w] = v820obus[temp_w*1 +:temp_w];
assign v820ibus[data_w*1 +:data_w] = c371obus[data_w*2 +:data_w];
assign c371ibus[temp_w*3 +:temp_w] = v876obus[temp_w*1 +:temp_w];
assign v876ibus[data_w*1 +:data_w] = c371obus[data_w*3 +:data_w];
assign c371ibus[temp_w*4 +:temp_w] = v1523obus[temp_w*1 +:temp_w];
assign v1523ibus[data_w*1 +:data_w] = c371obus[data_w*4 +:data_w];
assign c371ibus[temp_w*5 +:temp_w] = v1619obus[temp_w*0 +:temp_w];
assign v1619ibus[data_w*0 +:data_w] = c371obus[data_w*5 +:data_w];
assign c372ibus[temp_w*0 +:temp_w] = v49obus[temp_w*0 +:temp_w];
assign v49ibus[data_w*0 +:data_w] = c372obus[data_w*0 +:data_w];
assign c372ibus[temp_w*1 +:temp_w] = v227obus[temp_w*1 +:temp_w];
assign v227ibus[data_w*1 +:data_w] = c372obus[data_w*1 +:data_w];
assign c372ibus[temp_w*2 +:temp_w] = v821obus[temp_w*1 +:temp_w];
assign v821ibus[data_w*1 +:data_w] = c372obus[data_w*2 +:data_w];
assign c372ibus[temp_w*3 +:temp_w] = v877obus[temp_w*1 +:temp_w];
assign v877ibus[data_w*1 +:data_w] = c372obus[data_w*3 +:data_w];
assign c372ibus[temp_w*4 +:temp_w] = v1524obus[temp_w*1 +:temp_w];
assign v1524ibus[data_w*1 +:data_w] = c372obus[data_w*4 +:data_w];
assign c372ibus[temp_w*5 +:temp_w] = v1620obus[temp_w*0 +:temp_w];
assign v1620ibus[data_w*0 +:data_w] = c372obus[data_w*5 +:data_w];
assign c373ibus[temp_w*0 +:temp_w] = v50obus[temp_w*0 +:temp_w];
assign v50ibus[data_w*0 +:data_w] = c373obus[data_w*0 +:data_w];
assign c373ibus[temp_w*1 +:temp_w] = v228obus[temp_w*1 +:temp_w];
assign v228ibus[data_w*1 +:data_w] = c373obus[data_w*1 +:data_w];
assign c373ibus[temp_w*2 +:temp_w] = v822obus[temp_w*1 +:temp_w];
assign v822ibus[data_w*1 +:data_w] = c373obus[data_w*2 +:data_w];
assign c373ibus[temp_w*3 +:temp_w] = v878obus[temp_w*1 +:temp_w];
assign v878ibus[data_w*1 +:data_w] = c373obus[data_w*3 +:data_w];
assign c373ibus[temp_w*4 +:temp_w] = v1525obus[temp_w*1 +:temp_w];
assign v1525ibus[data_w*1 +:data_w] = c373obus[data_w*4 +:data_w];
assign c373ibus[temp_w*5 +:temp_w] = v1621obus[temp_w*0 +:temp_w];
assign v1621ibus[data_w*0 +:data_w] = c373obus[data_w*5 +:data_w];
assign c374ibus[temp_w*0 +:temp_w] = v51obus[temp_w*0 +:temp_w];
assign v51ibus[data_w*0 +:data_w] = c374obus[data_w*0 +:data_w];
assign c374ibus[temp_w*1 +:temp_w] = v229obus[temp_w*1 +:temp_w];
assign v229ibus[data_w*1 +:data_w] = c374obus[data_w*1 +:data_w];
assign c374ibus[temp_w*2 +:temp_w] = v823obus[temp_w*1 +:temp_w];
assign v823ibus[data_w*1 +:data_w] = c374obus[data_w*2 +:data_w];
assign c374ibus[temp_w*3 +:temp_w] = v879obus[temp_w*1 +:temp_w];
assign v879ibus[data_w*1 +:data_w] = c374obus[data_w*3 +:data_w];
assign c374ibus[temp_w*4 +:temp_w] = v1526obus[temp_w*1 +:temp_w];
assign v1526ibus[data_w*1 +:data_w] = c374obus[data_w*4 +:data_w];
assign c374ibus[temp_w*5 +:temp_w] = v1622obus[temp_w*0 +:temp_w];
assign v1622ibus[data_w*0 +:data_w] = c374obus[data_w*5 +:data_w];
assign c375ibus[temp_w*0 +:temp_w] = v52obus[temp_w*0 +:temp_w];
assign v52ibus[data_w*0 +:data_w] = c375obus[data_w*0 +:data_w];
assign c375ibus[temp_w*1 +:temp_w] = v230obus[temp_w*1 +:temp_w];
assign v230ibus[data_w*1 +:data_w] = c375obus[data_w*1 +:data_w];
assign c375ibus[temp_w*2 +:temp_w] = v824obus[temp_w*1 +:temp_w];
assign v824ibus[data_w*1 +:data_w] = c375obus[data_w*2 +:data_w];
assign c375ibus[temp_w*3 +:temp_w] = v880obus[temp_w*1 +:temp_w];
assign v880ibus[data_w*1 +:data_w] = c375obus[data_w*3 +:data_w];
assign c375ibus[temp_w*4 +:temp_w] = v1527obus[temp_w*1 +:temp_w];
assign v1527ibus[data_w*1 +:data_w] = c375obus[data_w*4 +:data_w];
assign c375ibus[temp_w*5 +:temp_w] = v1623obus[temp_w*0 +:temp_w];
assign v1623ibus[data_w*0 +:data_w] = c375obus[data_w*5 +:data_w];
assign c376ibus[temp_w*0 +:temp_w] = v53obus[temp_w*0 +:temp_w];
assign v53ibus[data_w*0 +:data_w] = c376obus[data_w*0 +:data_w];
assign c376ibus[temp_w*1 +:temp_w] = v231obus[temp_w*1 +:temp_w];
assign v231ibus[data_w*1 +:data_w] = c376obus[data_w*1 +:data_w];
assign c376ibus[temp_w*2 +:temp_w] = v825obus[temp_w*1 +:temp_w];
assign v825ibus[data_w*1 +:data_w] = c376obus[data_w*2 +:data_w];
assign c376ibus[temp_w*3 +:temp_w] = v881obus[temp_w*1 +:temp_w];
assign v881ibus[data_w*1 +:data_w] = c376obus[data_w*3 +:data_w];
assign c376ibus[temp_w*4 +:temp_w] = v1528obus[temp_w*1 +:temp_w];
assign v1528ibus[data_w*1 +:data_w] = c376obus[data_w*4 +:data_w];
assign c376ibus[temp_w*5 +:temp_w] = v1624obus[temp_w*0 +:temp_w];
assign v1624ibus[data_w*0 +:data_w] = c376obus[data_w*5 +:data_w];
assign c377ibus[temp_w*0 +:temp_w] = v54obus[temp_w*0 +:temp_w];
assign v54ibus[data_w*0 +:data_w] = c377obus[data_w*0 +:data_w];
assign c377ibus[temp_w*1 +:temp_w] = v232obus[temp_w*1 +:temp_w];
assign v232ibus[data_w*1 +:data_w] = c377obus[data_w*1 +:data_w];
assign c377ibus[temp_w*2 +:temp_w] = v826obus[temp_w*1 +:temp_w];
assign v826ibus[data_w*1 +:data_w] = c377obus[data_w*2 +:data_w];
assign c377ibus[temp_w*3 +:temp_w] = v882obus[temp_w*1 +:temp_w];
assign v882ibus[data_w*1 +:data_w] = c377obus[data_w*3 +:data_w];
assign c377ibus[temp_w*4 +:temp_w] = v1529obus[temp_w*1 +:temp_w];
assign v1529ibus[data_w*1 +:data_w] = c377obus[data_w*4 +:data_w];
assign c377ibus[temp_w*5 +:temp_w] = v1625obus[temp_w*0 +:temp_w];
assign v1625ibus[data_w*0 +:data_w] = c377obus[data_w*5 +:data_w];
assign c378ibus[temp_w*0 +:temp_w] = v55obus[temp_w*0 +:temp_w];
assign v55ibus[data_w*0 +:data_w] = c378obus[data_w*0 +:data_w];
assign c378ibus[temp_w*1 +:temp_w] = v233obus[temp_w*1 +:temp_w];
assign v233ibus[data_w*1 +:data_w] = c378obus[data_w*1 +:data_w];
assign c378ibus[temp_w*2 +:temp_w] = v827obus[temp_w*1 +:temp_w];
assign v827ibus[data_w*1 +:data_w] = c378obus[data_w*2 +:data_w];
assign c378ibus[temp_w*3 +:temp_w] = v883obus[temp_w*1 +:temp_w];
assign v883ibus[data_w*1 +:data_w] = c378obus[data_w*3 +:data_w];
assign c378ibus[temp_w*4 +:temp_w] = v1530obus[temp_w*1 +:temp_w];
assign v1530ibus[data_w*1 +:data_w] = c378obus[data_w*4 +:data_w];
assign c378ibus[temp_w*5 +:temp_w] = v1626obus[temp_w*0 +:temp_w];
assign v1626ibus[data_w*0 +:data_w] = c378obus[data_w*5 +:data_w];
assign c379ibus[temp_w*0 +:temp_w] = v56obus[temp_w*0 +:temp_w];
assign v56ibus[data_w*0 +:data_w] = c379obus[data_w*0 +:data_w];
assign c379ibus[temp_w*1 +:temp_w] = v234obus[temp_w*1 +:temp_w];
assign v234ibus[data_w*1 +:data_w] = c379obus[data_w*1 +:data_w];
assign c379ibus[temp_w*2 +:temp_w] = v828obus[temp_w*1 +:temp_w];
assign v828ibus[data_w*1 +:data_w] = c379obus[data_w*2 +:data_w];
assign c379ibus[temp_w*3 +:temp_w] = v884obus[temp_w*1 +:temp_w];
assign v884ibus[data_w*1 +:data_w] = c379obus[data_w*3 +:data_w];
assign c379ibus[temp_w*4 +:temp_w] = v1531obus[temp_w*1 +:temp_w];
assign v1531ibus[data_w*1 +:data_w] = c379obus[data_w*4 +:data_w];
assign c379ibus[temp_w*5 +:temp_w] = v1627obus[temp_w*0 +:temp_w];
assign v1627ibus[data_w*0 +:data_w] = c379obus[data_w*5 +:data_w];
assign c380ibus[temp_w*0 +:temp_w] = v57obus[temp_w*0 +:temp_w];
assign v57ibus[data_w*0 +:data_w] = c380obus[data_w*0 +:data_w];
assign c380ibus[temp_w*1 +:temp_w] = v235obus[temp_w*1 +:temp_w];
assign v235ibus[data_w*1 +:data_w] = c380obus[data_w*1 +:data_w];
assign c380ibus[temp_w*2 +:temp_w] = v829obus[temp_w*1 +:temp_w];
assign v829ibus[data_w*1 +:data_w] = c380obus[data_w*2 +:data_w];
assign c380ibus[temp_w*3 +:temp_w] = v885obus[temp_w*1 +:temp_w];
assign v885ibus[data_w*1 +:data_w] = c380obus[data_w*3 +:data_w];
assign c380ibus[temp_w*4 +:temp_w] = v1532obus[temp_w*1 +:temp_w];
assign v1532ibus[data_w*1 +:data_w] = c380obus[data_w*4 +:data_w];
assign c380ibus[temp_w*5 +:temp_w] = v1628obus[temp_w*0 +:temp_w];
assign v1628ibus[data_w*0 +:data_w] = c380obus[data_w*5 +:data_w];
assign c381ibus[temp_w*0 +:temp_w] = v58obus[temp_w*0 +:temp_w];
assign v58ibus[data_w*0 +:data_w] = c381obus[data_w*0 +:data_w];
assign c381ibus[temp_w*1 +:temp_w] = v236obus[temp_w*1 +:temp_w];
assign v236ibus[data_w*1 +:data_w] = c381obus[data_w*1 +:data_w];
assign c381ibus[temp_w*2 +:temp_w] = v830obus[temp_w*1 +:temp_w];
assign v830ibus[data_w*1 +:data_w] = c381obus[data_w*2 +:data_w];
assign c381ibus[temp_w*3 +:temp_w] = v886obus[temp_w*1 +:temp_w];
assign v886ibus[data_w*1 +:data_w] = c381obus[data_w*3 +:data_w];
assign c381ibus[temp_w*4 +:temp_w] = v1533obus[temp_w*1 +:temp_w];
assign v1533ibus[data_w*1 +:data_w] = c381obus[data_w*4 +:data_w];
assign c381ibus[temp_w*5 +:temp_w] = v1629obus[temp_w*0 +:temp_w];
assign v1629ibus[data_w*0 +:data_w] = c381obus[data_w*5 +:data_w];
assign c382ibus[temp_w*0 +:temp_w] = v59obus[temp_w*0 +:temp_w];
assign v59ibus[data_w*0 +:data_w] = c382obus[data_w*0 +:data_w];
assign c382ibus[temp_w*1 +:temp_w] = v237obus[temp_w*1 +:temp_w];
assign v237ibus[data_w*1 +:data_w] = c382obus[data_w*1 +:data_w];
assign c382ibus[temp_w*2 +:temp_w] = v831obus[temp_w*1 +:temp_w];
assign v831ibus[data_w*1 +:data_w] = c382obus[data_w*2 +:data_w];
assign c382ibus[temp_w*3 +:temp_w] = v887obus[temp_w*1 +:temp_w];
assign v887ibus[data_w*1 +:data_w] = c382obus[data_w*3 +:data_w];
assign c382ibus[temp_w*4 +:temp_w] = v1534obus[temp_w*1 +:temp_w];
assign v1534ibus[data_w*1 +:data_w] = c382obus[data_w*4 +:data_w];
assign c382ibus[temp_w*5 +:temp_w] = v1630obus[temp_w*0 +:temp_w];
assign v1630ibus[data_w*0 +:data_w] = c382obus[data_w*5 +:data_w];
assign c383ibus[temp_w*0 +:temp_w] = v60obus[temp_w*0 +:temp_w];
assign v60ibus[data_w*0 +:data_w] = c383obus[data_w*0 +:data_w];
assign c383ibus[temp_w*1 +:temp_w] = v238obus[temp_w*1 +:temp_w];
assign v238ibus[data_w*1 +:data_w] = c383obus[data_w*1 +:data_w];
assign c383ibus[temp_w*2 +:temp_w] = v832obus[temp_w*1 +:temp_w];
assign v832ibus[data_w*1 +:data_w] = c383obus[data_w*2 +:data_w];
assign c383ibus[temp_w*3 +:temp_w] = v888obus[temp_w*1 +:temp_w];
assign v888ibus[data_w*1 +:data_w] = c383obus[data_w*3 +:data_w];
assign c383ibus[temp_w*4 +:temp_w] = v1535obus[temp_w*1 +:temp_w];
assign v1535ibus[data_w*1 +:data_w] = c383obus[data_w*4 +:data_w];
assign c383ibus[temp_w*5 +:temp_w] = v1631obus[temp_w*0 +:temp_w];
assign v1631ibus[data_w*0 +:data_w] = c383obus[data_w*5 +:data_w];
assign c384ibus[temp_w*0 +:temp_w] = v231obus[temp_w*2 +:temp_w];
assign v231ibus[data_w*2 +:data_w] = c384obus[data_w*0 +:data_w];
assign c384ibus[temp_w*1 +:temp_w] = v660obus[temp_w*1 +:temp_w];
assign v660ibus[data_w*1 +:data_w] = c384obus[data_w*1 +:data_w];
assign c384ibus[temp_w*2 +:temp_w] = v905obus[temp_w*2 +:temp_w];
assign v905ibus[data_w*2 +:data_w] = c384obus[data_w*2 +:data_w];
assign c384ibus[temp_w*3 +:temp_w] = v1032obus[temp_w*0 +:temp_w];
assign v1032ibus[data_w*0 +:data_w] = c384obus[data_w*3 +:data_w];
assign c384ibus[temp_w*4 +:temp_w] = v1536obus[temp_w*1 +:temp_w];
assign v1536ibus[data_w*1 +:data_w] = c384obus[data_w*4 +:data_w];
assign c384ibus[temp_w*5 +:temp_w] = v1632obus[temp_w*0 +:temp_w];
assign v1632ibus[data_w*0 +:data_w] = c384obus[data_w*5 +:data_w];
assign c385ibus[temp_w*0 +:temp_w] = v232obus[temp_w*2 +:temp_w];
assign v232ibus[data_w*2 +:data_w] = c385obus[data_w*0 +:data_w];
assign c385ibus[temp_w*1 +:temp_w] = v661obus[temp_w*1 +:temp_w];
assign v661ibus[data_w*1 +:data_w] = c385obus[data_w*1 +:data_w];
assign c385ibus[temp_w*2 +:temp_w] = v906obus[temp_w*2 +:temp_w];
assign v906ibus[data_w*2 +:data_w] = c385obus[data_w*2 +:data_w];
assign c385ibus[temp_w*3 +:temp_w] = v1033obus[temp_w*0 +:temp_w];
assign v1033ibus[data_w*0 +:data_w] = c385obus[data_w*3 +:data_w];
assign c385ibus[temp_w*4 +:temp_w] = v1537obus[temp_w*1 +:temp_w];
assign v1537ibus[data_w*1 +:data_w] = c385obus[data_w*4 +:data_w];
assign c385ibus[temp_w*5 +:temp_w] = v1633obus[temp_w*0 +:temp_w];
assign v1633ibus[data_w*0 +:data_w] = c385obus[data_w*5 +:data_w];
assign c386ibus[temp_w*0 +:temp_w] = v233obus[temp_w*2 +:temp_w];
assign v233ibus[data_w*2 +:data_w] = c386obus[data_w*0 +:data_w];
assign c386ibus[temp_w*1 +:temp_w] = v662obus[temp_w*1 +:temp_w];
assign v662ibus[data_w*1 +:data_w] = c386obus[data_w*1 +:data_w];
assign c386ibus[temp_w*2 +:temp_w] = v907obus[temp_w*2 +:temp_w];
assign v907ibus[data_w*2 +:data_w] = c386obus[data_w*2 +:data_w];
assign c386ibus[temp_w*3 +:temp_w] = v1034obus[temp_w*0 +:temp_w];
assign v1034ibus[data_w*0 +:data_w] = c386obus[data_w*3 +:data_w];
assign c386ibus[temp_w*4 +:temp_w] = v1538obus[temp_w*1 +:temp_w];
assign v1538ibus[data_w*1 +:data_w] = c386obus[data_w*4 +:data_w];
assign c386ibus[temp_w*5 +:temp_w] = v1634obus[temp_w*0 +:temp_w];
assign v1634ibus[data_w*0 +:data_w] = c386obus[data_w*5 +:data_w];
assign c387ibus[temp_w*0 +:temp_w] = v234obus[temp_w*2 +:temp_w];
assign v234ibus[data_w*2 +:data_w] = c387obus[data_w*0 +:data_w];
assign c387ibus[temp_w*1 +:temp_w] = v663obus[temp_w*1 +:temp_w];
assign v663ibus[data_w*1 +:data_w] = c387obus[data_w*1 +:data_w];
assign c387ibus[temp_w*2 +:temp_w] = v908obus[temp_w*2 +:temp_w];
assign v908ibus[data_w*2 +:data_w] = c387obus[data_w*2 +:data_w];
assign c387ibus[temp_w*3 +:temp_w] = v1035obus[temp_w*0 +:temp_w];
assign v1035ibus[data_w*0 +:data_w] = c387obus[data_w*3 +:data_w];
assign c387ibus[temp_w*4 +:temp_w] = v1539obus[temp_w*1 +:temp_w];
assign v1539ibus[data_w*1 +:data_w] = c387obus[data_w*4 +:data_w];
assign c387ibus[temp_w*5 +:temp_w] = v1635obus[temp_w*0 +:temp_w];
assign v1635ibus[data_w*0 +:data_w] = c387obus[data_w*5 +:data_w];
assign c388ibus[temp_w*0 +:temp_w] = v235obus[temp_w*2 +:temp_w];
assign v235ibus[data_w*2 +:data_w] = c388obus[data_w*0 +:data_w];
assign c388ibus[temp_w*1 +:temp_w] = v664obus[temp_w*1 +:temp_w];
assign v664ibus[data_w*1 +:data_w] = c388obus[data_w*1 +:data_w];
assign c388ibus[temp_w*2 +:temp_w] = v909obus[temp_w*2 +:temp_w];
assign v909ibus[data_w*2 +:data_w] = c388obus[data_w*2 +:data_w];
assign c388ibus[temp_w*3 +:temp_w] = v1036obus[temp_w*0 +:temp_w];
assign v1036ibus[data_w*0 +:data_w] = c388obus[data_w*3 +:data_w];
assign c388ibus[temp_w*4 +:temp_w] = v1540obus[temp_w*1 +:temp_w];
assign v1540ibus[data_w*1 +:data_w] = c388obus[data_w*4 +:data_w];
assign c388ibus[temp_w*5 +:temp_w] = v1636obus[temp_w*0 +:temp_w];
assign v1636ibus[data_w*0 +:data_w] = c388obus[data_w*5 +:data_w];
assign c389ibus[temp_w*0 +:temp_w] = v236obus[temp_w*2 +:temp_w];
assign v236ibus[data_w*2 +:data_w] = c389obus[data_w*0 +:data_w];
assign c389ibus[temp_w*1 +:temp_w] = v665obus[temp_w*1 +:temp_w];
assign v665ibus[data_w*1 +:data_w] = c389obus[data_w*1 +:data_w];
assign c389ibus[temp_w*2 +:temp_w] = v910obus[temp_w*2 +:temp_w];
assign v910ibus[data_w*2 +:data_w] = c389obus[data_w*2 +:data_w];
assign c389ibus[temp_w*3 +:temp_w] = v1037obus[temp_w*0 +:temp_w];
assign v1037ibus[data_w*0 +:data_w] = c389obus[data_w*3 +:data_w];
assign c389ibus[temp_w*4 +:temp_w] = v1541obus[temp_w*1 +:temp_w];
assign v1541ibus[data_w*1 +:data_w] = c389obus[data_w*4 +:data_w];
assign c389ibus[temp_w*5 +:temp_w] = v1637obus[temp_w*0 +:temp_w];
assign v1637ibus[data_w*0 +:data_w] = c389obus[data_w*5 +:data_w];
assign c390ibus[temp_w*0 +:temp_w] = v237obus[temp_w*2 +:temp_w];
assign v237ibus[data_w*2 +:data_w] = c390obus[data_w*0 +:data_w];
assign c390ibus[temp_w*1 +:temp_w] = v666obus[temp_w*1 +:temp_w];
assign v666ibus[data_w*1 +:data_w] = c390obus[data_w*1 +:data_w];
assign c390ibus[temp_w*2 +:temp_w] = v911obus[temp_w*2 +:temp_w];
assign v911ibus[data_w*2 +:data_w] = c390obus[data_w*2 +:data_w];
assign c390ibus[temp_w*3 +:temp_w] = v1038obus[temp_w*0 +:temp_w];
assign v1038ibus[data_w*0 +:data_w] = c390obus[data_w*3 +:data_w];
assign c390ibus[temp_w*4 +:temp_w] = v1542obus[temp_w*1 +:temp_w];
assign v1542ibus[data_w*1 +:data_w] = c390obus[data_w*4 +:data_w];
assign c390ibus[temp_w*5 +:temp_w] = v1638obus[temp_w*0 +:temp_w];
assign v1638ibus[data_w*0 +:data_w] = c390obus[data_w*5 +:data_w];
assign c391ibus[temp_w*0 +:temp_w] = v238obus[temp_w*2 +:temp_w];
assign v238ibus[data_w*2 +:data_w] = c391obus[data_w*0 +:data_w];
assign c391ibus[temp_w*1 +:temp_w] = v667obus[temp_w*1 +:temp_w];
assign v667ibus[data_w*1 +:data_w] = c391obus[data_w*1 +:data_w];
assign c391ibus[temp_w*2 +:temp_w] = v912obus[temp_w*2 +:temp_w];
assign v912ibus[data_w*2 +:data_w] = c391obus[data_w*2 +:data_w];
assign c391ibus[temp_w*3 +:temp_w] = v1039obus[temp_w*0 +:temp_w];
assign v1039ibus[data_w*0 +:data_w] = c391obus[data_w*3 +:data_w];
assign c391ibus[temp_w*4 +:temp_w] = v1543obus[temp_w*1 +:temp_w];
assign v1543ibus[data_w*1 +:data_w] = c391obus[data_w*4 +:data_w];
assign c391ibus[temp_w*5 +:temp_w] = v1639obus[temp_w*0 +:temp_w];
assign v1639ibus[data_w*0 +:data_w] = c391obus[data_w*5 +:data_w];
assign c392ibus[temp_w*0 +:temp_w] = v239obus[temp_w*2 +:temp_w];
assign v239ibus[data_w*2 +:data_w] = c392obus[data_w*0 +:data_w];
assign c392ibus[temp_w*1 +:temp_w] = v668obus[temp_w*1 +:temp_w];
assign v668ibus[data_w*1 +:data_w] = c392obus[data_w*1 +:data_w];
assign c392ibus[temp_w*2 +:temp_w] = v913obus[temp_w*2 +:temp_w];
assign v913ibus[data_w*2 +:data_w] = c392obus[data_w*2 +:data_w];
assign c392ibus[temp_w*3 +:temp_w] = v1040obus[temp_w*0 +:temp_w];
assign v1040ibus[data_w*0 +:data_w] = c392obus[data_w*3 +:data_w];
assign c392ibus[temp_w*4 +:temp_w] = v1544obus[temp_w*1 +:temp_w];
assign v1544ibus[data_w*1 +:data_w] = c392obus[data_w*4 +:data_w];
assign c392ibus[temp_w*5 +:temp_w] = v1640obus[temp_w*0 +:temp_w];
assign v1640ibus[data_w*0 +:data_w] = c392obus[data_w*5 +:data_w];
assign c393ibus[temp_w*0 +:temp_w] = v240obus[temp_w*2 +:temp_w];
assign v240ibus[data_w*2 +:data_w] = c393obus[data_w*0 +:data_w];
assign c393ibus[temp_w*1 +:temp_w] = v669obus[temp_w*1 +:temp_w];
assign v669ibus[data_w*1 +:data_w] = c393obus[data_w*1 +:data_w];
assign c393ibus[temp_w*2 +:temp_w] = v914obus[temp_w*2 +:temp_w];
assign v914ibus[data_w*2 +:data_w] = c393obus[data_w*2 +:data_w];
assign c393ibus[temp_w*3 +:temp_w] = v1041obus[temp_w*0 +:temp_w];
assign v1041ibus[data_w*0 +:data_w] = c393obus[data_w*3 +:data_w];
assign c393ibus[temp_w*4 +:temp_w] = v1545obus[temp_w*1 +:temp_w];
assign v1545ibus[data_w*1 +:data_w] = c393obus[data_w*4 +:data_w];
assign c393ibus[temp_w*5 +:temp_w] = v1641obus[temp_w*0 +:temp_w];
assign v1641ibus[data_w*0 +:data_w] = c393obus[data_w*5 +:data_w];
assign c394ibus[temp_w*0 +:temp_w] = v241obus[temp_w*2 +:temp_w];
assign v241ibus[data_w*2 +:data_w] = c394obus[data_w*0 +:data_w];
assign c394ibus[temp_w*1 +:temp_w] = v670obus[temp_w*1 +:temp_w];
assign v670ibus[data_w*1 +:data_w] = c394obus[data_w*1 +:data_w];
assign c394ibus[temp_w*2 +:temp_w] = v915obus[temp_w*2 +:temp_w];
assign v915ibus[data_w*2 +:data_w] = c394obus[data_w*2 +:data_w];
assign c394ibus[temp_w*3 +:temp_w] = v1042obus[temp_w*0 +:temp_w];
assign v1042ibus[data_w*0 +:data_w] = c394obus[data_w*3 +:data_w];
assign c394ibus[temp_w*4 +:temp_w] = v1546obus[temp_w*1 +:temp_w];
assign v1546ibus[data_w*1 +:data_w] = c394obus[data_w*4 +:data_w];
assign c394ibus[temp_w*5 +:temp_w] = v1642obus[temp_w*0 +:temp_w];
assign v1642ibus[data_w*0 +:data_w] = c394obus[data_w*5 +:data_w];
assign c395ibus[temp_w*0 +:temp_w] = v242obus[temp_w*2 +:temp_w];
assign v242ibus[data_w*2 +:data_w] = c395obus[data_w*0 +:data_w];
assign c395ibus[temp_w*1 +:temp_w] = v671obus[temp_w*1 +:temp_w];
assign v671ibus[data_w*1 +:data_w] = c395obus[data_w*1 +:data_w];
assign c395ibus[temp_w*2 +:temp_w] = v916obus[temp_w*2 +:temp_w];
assign v916ibus[data_w*2 +:data_w] = c395obus[data_w*2 +:data_w];
assign c395ibus[temp_w*3 +:temp_w] = v1043obus[temp_w*0 +:temp_w];
assign v1043ibus[data_w*0 +:data_w] = c395obus[data_w*3 +:data_w];
assign c395ibus[temp_w*4 +:temp_w] = v1547obus[temp_w*1 +:temp_w];
assign v1547ibus[data_w*1 +:data_w] = c395obus[data_w*4 +:data_w];
assign c395ibus[temp_w*5 +:temp_w] = v1643obus[temp_w*0 +:temp_w];
assign v1643ibus[data_w*0 +:data_w] = c395obus[data_w*5 +:data_w];
assign c396ibus[temp_w*0 +:temp_w] = v243obus[temp_w*2 +:temp_w];
assign v243ibus[data_w*2 +:data_w] = c396obus[data_w*0 +:data_w];
assign c396ibus[temp_w*1 +:temp_w] = v576obus[temp_w*1 +:temp_w];
assign v576ibus[data_w*1 +:data_w] = c396obus[data_w*1 +:data_w];
assign c396ibus[temp_w*2 +:temp_w] = v917obus[temp_w*2 +:temp_w];
assign v917ibus[data_w*2 +:data_w] = c396obus[data_w*2 +:data_w];
assign c396ibus[temp_w*3 +:temp_w] = v1044obus[temp_w*0 +:temp_w];
assign v1044ibus[data_w*0 +:data_w] = c396obus[data_w*3 +:data_w];
assign c396ibus[temp_w*4 +:temp_w] = v1548obus[temp_w*1 +:temp_w];
assign v1548ibus[data_w*1 +:data_w] = c396obus[data_w*4 +:data_w];
assign c396ibus[temp_w*5 +:temp_w] = v1644obus[temp_w*0 +:temp_w];
assign v1644ibus[data_w*0 +:data_w] = c396obus[data_w*5 +:data_w];
assign c397ibus[temp_w*0 +:temp_w] = v244obus[temp_w*2 +:temp_w];
assign v244ibus[data_w*2 +:data_w] = c397obus[data_w*0 +:data_w];
assign c397ibus[temp_w*1 +:temp_w] = v577obus[temp_w*1 +:temp_w];
assign v577ibus[data_w*1 +:data_w] = c397obus[data_w*1 +:data_w];
assign c397ibus[temp_w*2 +:temp_w] = v918obus[temp_w*2 +:temp_w];
assign v918ibus[data_w*2 +:data_w] = c397obus[data_w*2 +:data_w];
assign c397ibus[temp_w*3 +:temp_w] = v1045obus[temp_w*0 +:temp_w];
assign v1045ibus[data_w*0 +:data_w] = c397obus[data_w*3 +:data_w];
assign c397ibus[temp_w*4 +:temp_w] = v1549obus[temp_w*1 +:temp_w];
assign v1549ibus[data_w*1 +:data_w] = c397obus[data_w*4 +:data_w];
assign c397ibus[temp_w*5 +:temp_w] = v1645obus[temp_w*0 +:temp_w];
assign v1645ibus[data_w*0 +:data_w] = c397obus[data_w*5 +:data_w];
assign c398ibus[temp_w*0 +:temp_w] = v245obus[temp_w*2 +:temp_w];
assign v245ibus[data_w*2 +:data_w] = c398obus[data_w*0 +:data_w];
assign c398ibus[temp_w*1 +:temp_w] = v578obus[temp_w*1 +:temp_w];
assign v578ibus[data_w*1 +:data_w] = c398obus[data_w*1 +:data_w];
assign c398ibus[temp_w*2 +:temp_w] = v919obus[temp_w*2 +:temp_w];
assign v919ibus[data_w*2 +:data_w] = c398obus[data_w*2 +:data_w];
assign c398ibus[temp_w*3 +:temp_w] = v1046obus[temp_w*0 +:temp_w];
assign v1046ibus[data_w*0 +:data_w] = c398obus[data_w*3 +:data_w];
assign c398ibus[temp_w*4 +:temp_w] = v1550obus[temp_w*1 +:temp_w];
assign v1550ibus[data_w*1 +:data_w] = c398obus[data_w*4 +:data_w];
assign c398ibus[temp_w*5 +:temp_w] = v1646obus[temp_w*0 +:temp_w];
assign v1646ibus[data_w*0 +:data_w] = c398obus[data_w*5 +:data_w];
assign c399ibus[temp_w*0 +:temp_w] = v246obus[temp_w*2 +:temp_w];
assign v246ibus[data_w*2 +:data_w] = c399obus[data_w*0 +:data_w];
assign c399ibus[temp_w*1 +:temp_w] = v579obus[temp_w*1 +:temp_w];
assign v579ibus[data_w*1 +:data_w] = c399obus[data_w*1 +:data_w];
assign c399ibus[temp_w*2 +:temp_w] = v920obus[temp_w*2 +:temp_w];
assign v920ibus[data_w*2 +:data_w] = c399obus[data_w*2 +:data_w];
assign c399ibus[temp_w*3 +:temp_w] = v1047obus[temp_w*0 +:temp_w];
assign v1047ibus[data_w*0 +:data_w] = c399obus[data_w*3 +:data_w];
assign c399ibus[temp_w*4 +:temp_w] = v1551obus[temp_w*1 +:temp_w];
assign v1551ibus[data_w*1 +:data_w] = c399obus[data_w*4 +:data_w];
assign c399ibus[temp_w*5 +:temp_w] = v1647obus[temp_w*0 +:temp_w];
assign v1647ibus[data_w*0 +:data_w] = c399obus[data_w*5 +:data_w];
assign c400ibus[temp_w*0 +:temp_w] = v247obus[temp_w*2 +:temp_w];
assign v247ibus[data_w*2 +:data_w] = c400obus[data_w*0 +:data_w];
assign c400ibus[temp_w*1 +:temp_w] = v580obus[temp_w*1 +:temp_w];
assign v580ibus[data_w*1 +:data_w] = c400obus[data_w*1 +:data_w];
assign c400ibus[temp_w*2 +:temp_w] = v921obus[temp_w*2 +:temp_w];
assign v921ibus[data_w*2 +:data_w] = c400obus[data_w*2 +:data_w];
assign c400ibus[temp_w*3 +:temp_w] = v1048obus[temp_w*0 +:temp_w];
assign v1048ibus[data_w*0 +:data_w] = c400obus[data_w*3 +:data_w];
assign c400ibus[temp_w*4 +:temp_w] = v1552obus[temp_w*1 +:temp_w];
assign v1552ibus[data_w*1 +:data_w] = c400obus[data_w*4 +:data_w];
assign c400ibus[temp_w*5 +:temp_w] = v1648obus[temp_w*0 +:temp_w];
assign v1648ibus[data_w*0 +:data_w] = c400obus[data_w*5 +:data_w];
assign c401ibus[temp_w*0 +:temp_w] = v248obus[temp_w*2 +:temp_w];
assign v248ibus[data_w*2 +:data_w] = c401obus[data_w*0 +:data_w];
assign c401ibus[temp_w*1 +:temp_w] = v581obus[temp_w*1 +:temp_w];
assign v581ibus[data_w*1 +:data_w] = c401obus[data_w*1 +:data_w];
assign c401ibus[temp_w*2 +:temp_w] = v922obus[temp_w*2 +:temp_w];
assign v922ibus[data_w*2 +:data_w] = c401obus[data_w*2 +:data_w];
assign c401ibus[temp_w*3 +:temp_w] = v1049obus[temp_w*0 +:temp_w];
assign v1049ibus[data_w*0 +:data_w] = c401obus[data_w*3 +:data_w];
assign c401ibus[temp_w*4 +:temp_w] = v1553obus[temp_w*1 +:temp_w];
assign v1553ibus[data_w*1 +:data_w] = c401obus[data_w*4 +:data_w];
assign c401ibus[temp_w*5 +:temp_w] = v1649obus[temp_w*0 +:temp_w];
assign v1649ibus[data_w*0 +:data_w] = c401obus[data_w*5 +:data_w];
assign c402ibus[temp_w*0 +:temp_w] = v249obus[temp_w*2 +:temp_w];
assign v249ibus[data_w*2 +:data_w] = c402obus[data_w*0 +:data_w];
assign c402ibus[temp_w*1 +:temp_w] = v582obus[temp_w*1 +:temp_w];
assign v582ibus[data_w*1 +:data_w] = c402obus[data_w*1 +:data_w];
assign c402ibus[temp_w*2 +:temp_w] = v923obus[temp_w*2 +:temp_w];
assign v923ibus[data_w*2 +:data_w] = c402obus[data_w*2 +:data_w];
assign c402ibus[temp_w*3 +:temp_w] = v1050obus[temp_w*0 +:temp_w];
assign v1050ibus[data_w*0 +:data_w] = c402obus[data_w*3 +:data_w];
assign c402ibus[temp_w*4 +:temp_w] = v1554obus[temp_w*1 +:temp_w];
assign v1554ibus[data_w*1 +:data_w] = c402obus[data_w*4 +:data_w];
assign c402ibus[temp_w*5 +:temp_w] = v1650obus[temp_w*0 +:temp_w];
assign v1650ibus[data_w*0 +:data_w] = c402obus[data_w*5 +:data_w];
assign c403ibus[temp_w*0 +:temp_w] = v250obus[temp_w*2 +:temp_w];
assign v250ibus[data_w*2 +:data_w] = c403obus[data_w*0 +:data_w];
assign c403ibus[temp_w*1 +:temp_w] = v583obus[temp_w*1 +:temp_w];
assign v583ibus[data_w*1 +:data_w] = c403obus[data_w*1 +:data_w];
assign c403ibus[temp_w*2 +:temp_w] = v924obus[temp_w*2 +:temp_w];
assign v924ibus[data_w*2 +:data_w] = c403obus[data_w*2 +:data_w];
assign c403ibus[temp_w*3 +:temp_w] = v1051obus[temp_w*0 +:temp_w];
assign v1051ibus[data_w*0 +:data_w] = c403obus[data_w*3 +:data_w];
assign c403ibus[temp_w*4 +:temp_w] = v1555obus[temp_w*1 +:temp_w];
assign v1555ibus[data_w*1 +:data_w] = c403obus[data_w*4 +:data_w];
assign c403ibus[temp_w*5 +:temp_w] = v1651obus[temp_w*0 +:temp_w];
assign v1651ibus[data_w*0 +:data_w] = c403obus[data_w*5 +:data_w];
assign c404ibus[temp_w*0 +:temp_w] = v251obus[temp_w*2 +:temp_w];
assign v251ibus[data_w*2 +:data_w] = c404obus[data_w*0 +:data_w];
assign c404ibus[temp_w*1 +:temp_w] = v584obus[temp_w*1 +:temp_w];
assign v584ibus[data_w*1 +:data_w] = c404obus[data_w*1 +:data_w];
assign c404ibus[temp_w*2 +:temp_w] = v925obus[temp_w*2 +:temp_w];
assign v925ibus[data_w*2 +:data_w] = c404obus[data_w*2 +:data_w];
assign c404ibus[temp_w*3 +:temp_w] = v1052obus[temp_w*0 +:temp_w];
assign v1052ibus[data_w*0 +:data_w] = c404obus[data_w*3 +:data_w];
assign c404ibus[temp_w*4 +:temp_w] = v1556obus[temp_w*1 +:temp_w];
assign v1556ibus[data_w*1 +:data_w] = c404obus[data_w*4 +:data_w];
assign c404ibus[temp_w*5 +:temp_w] = v1652obus[temp_w*0 +:temp_w];
assign v1652ibus[data_w*0 +:data_w] = c404obus[data_w*5 +:data_w];
assign c405ibus[temp_w*0 +:temp_w] = v252obus[temp_w*2 +:temp_w];
assign v252ibus[data_w*2 +:data_w] = c405obus[data_w*0 +:data_w];
assign c405ibus[temp_w*1 +:temp_w] = v585obus[temp_w*1 +:temp_w];
assign v585ibus[data_w*1 +:data_w] = c405obus[data_w*1 +:data_w];
assign c405ibus[temp_w*2 +:temp_w] = v926obus[temp_w*2 +:temp_w];
assign v926ibus[data_w*2 +:data_w] = c405obus[data_w*2 +:data_w];
assign c405ibus[temp_w*3 +:temp_w] = v1053obus[temp_w*0 +:temp_w];
assign v1053ibus[data_w*0 +:data_w] = c405obus[data_w*3 +:data_w];
assign c405ibus[temp_w*4 +:temp_w] = v1557obus[temp_w*1 +:temp_w];
assign v1557ibus[data_w*1 +:data_w] = c405obus[data_w*4 +:data_w];
assign c405ibus[temp_w*5 +:temp_w] = v1653obus[temp_w*0 +:temp_w];
assign v1653ibus[data_w*0 +:data_w] = c405obus[data_w*5 +:data_w];
assign c406ibus[temp_w*0 +:temp_w] = v253obus[temp_w*2 +:temp_w];
assign v253ibus[data_w*2 +:data_w] = c406obus[data_w*0 +:data_w];
assign c406ibus[temp_w*1 +:temp_w] = v586obus[temp_w*1 +:temp_w];
assign v586ibus[data_w*1 +:data_w] = c406obus[data_w*1 +:data_w];
assign c406ibus[temp_w*2 +:temp_w] = v927obus[temp_w*2 +:temp_w];
assign v927ibus[data_w*2 +:data_w] = c406obus[data_w*2 +:data_w];
assign c406ibus[temp_w*3 +:temp_w] = v1054obus[temp_w*0 +:temp_w];
assign v1054ibus[data_w*0 +:data_w] = c406obus[data_w*3 +:data_w];
assign c406ibus[temp_w*4 +:temp_w] = v1558obus[temp_w*1 +:temp_w];
assign v1558ibus[data_w*1 +:data_w] = c406obus[data_w*4 +:data_w];
assign c406ibus[temp_w*5 +:temp_w] = v1654obus[temp_w*0 +:temp_w];
assign v1654ibus[data_w*0 +:data_w] = c406obus[data_w*5 +:data_w];
assign c407ibus[temp_w*0 +:temp_w] = v254obus[temp_w*2 +:temp_w];
assign v254ibus[data_w*2 +:data_w] = c407obus[data_w*0 +:data_w];
assign c407ibus[temp_w*1 +:temp_w] = v587obus[temp_w*1 +:temp_w];
assign v587ibus[data_w*1 +:data_w] = c407obus[data_w*1 +:data_w];
assign c407ibus[temp_w*2 +:temp_w] = v928obus[temp_w*2 +:temp_w];
assign v928ibus[data_w*2 +:data_w] = c407obus[data_w*2 +:data_w];
assign c407ibus[temp_w*3 +:temp_w] = v1055obus[temp_w*0 +:temp_w];
assign v1055ibus[data_w*0 +:data_w] = c407obus[data_w*3 +:data_w];
assign c407ibus[temp_w*4 +:temp_w] = v1559obus[temp_w*1 +:temp_w];
assign v1559ibus[data_w*1 +:data_w] = c407obus[data_w*4 +:data_w];
assign c407ibus[temp_w*5 +:temp_w] = v1655obus[temp_w*0 +:temp_w];
assign v1655ibus[data_w*0 +:data_w] = c407obus[data_w*5 +:data_w];
assign c408ibus[temp_w*0 +:temp_w] = v255obus[temp_w*2 +:temp_w];
assign v255ibus[data_w*2 +:data_w] = c408obus[data_w*0 +:data_w];
assign c408ibus[temp_w*1 +:temp_w] = v588obus[temp_w*1 +:temp_w];
assign v588ibus[data_w*1 +:data_w] = c408obus[data_w*1 +:data_w];
assign c408ibus[temp_w*2 +:temp_w] = v929obus[temp_w*2 +:temp_w];
assign v929ibus[data_w*2 +:data_w] = c408obus[data_w*2 +:data_w];
assign c408ibus[temp_w*3 +:temp_w] = v960obus[temp_w*0 +:temp_w];
assign v960ibus[data_w*0 +:data_w] = c408obus[data_w*3 +:data_w];
assign c408ibus[temp_w*4 +:temp_w] = v1560obus[temp_w*1 +:temp_w];
assign v1560ibus[data_w*1 +:data_w] = c408obus[data_w*4 +:data_w];
assign c408ibus[temp_w*5 +:temp_w] = v1656obus[temp_w*0 +:temp_w];
assign v1656ibus[data_w*0 +:data_w] = c408obus[data_w*5 +:data_w];
assign c409ibus[temp_w*0 +:temp_w] = v256obus[temp_w*2 +:temp_w];
assign v256ibus[data_w*2 +:data_w] = c409obus[data_w*0 +:data_w];
assign c409ibus[temp_w*1 +:temp_w] = v589obus[temp_w*1 +:temp_w];
assign v589ibus[data_w*1 +:data_w] = c409obus[data_w*1 +:data_w];
assign c409ibus[temp_w*2 +:temp_w] = v930obus[temp_w*2 +:temp_w];
assign v930ibus[data_w*2 +:data_w] = c409obus[data_w*2 +:data_w];
assign c409ibus[temp_w*3 +:temp_w] = v961obus[temp_w*0 +:temp_w];
assign v961ibus[data_w*0 +:data_w] = c409obus[data_w*3 +:data_w];
assign c409ibus[temp_w*4 +:temp_w] = v1561obus[temp_w*1 +:temp_w];
assign v1561ibus[data_w*1 +:data_w] = c409obus[data_w*4 +:data_w];
assign c409ibus[temp_w*5 +:temp_w] = v1657obus[temp_w*0 +:temp_w];
assign v1657ibus[data_w*0 +:data_w] = c409obus[data_w*5 +:data_w];
assign c410ibus[temp_w*0 +:temp_w] = v257obus[temp_w*2 +:temp_w];
assign v257ibus[data_w*2 +:data_w] = c410obus[data_w*0 +:data_w];
assign c410ibus[temp_w*1 +:temp_w] = v590obus[temp_w*1 +:temp_w];
assign v590ibus[data_w*1 +:data_w] = c410obus[data_w*1 +:data_w];
assign c410ibus[temp_w*2 +:temp_w] = v931obus[temp_w*2 +:temp_w];
assign v931ibus[data_w*2 +:data_w] = c410obus[data_w*2 +:data_w];
assign c410ibus[temp_w*3 +:temp_w] = v962obus[temp_w*0 +:temp_w];
assign v962ibus[data_w*0 +:data_w] = c410obus[data_w*3 +:data_w];
assign c410ibus[temp_w*4 +:temp_w] = v1562obus[temp_w*1 +:temp_w];
assign v1562ibus[data_w*1 +:data_w] = c410obus[data_w*4 +:data_w];
assign c410ibus[temp_w*5 +:temp_w] = v1658obus[temp_w*0 +:temp_w];
assign v1658ibus[data_w*0 +:data_w] = c410obus[data_w*5 +:data_w];
assign c411ibus[temp_w*0 +:temp_w] = v258obus[temp_w*2 +:temp_w];
assign v258ibus[data_w*2 +:data_w] = c411obus[data_w*0 +:data_w];
assign c411ibus[temp_w*1 +:temp_w] = v591obus[temp_w*1 +:temp_w];
assign v591ibus[data_w*1 +:data_w] = c411obus[data_w*1 +:data_w];
assign c411ibus[temp_w*2 +:temp_w] = v932obus[temp_w*2 +:temp_w];
assign v932ibus[data_w*2 +:data_w] = c411obus[data_w*2 +:data_w];
assign c411ibus[temp_w*3 +:temp_w] = v963obus[temp_w*0 +:temp_w];
assign v963ibus[data_w*0 +:data_w] = c411obus[data_w*3 +:data_w];
assign c411ibus[temp_w*4 +:temp_w] = v1563obus[temp_w*1 +:temp_w];
assign v1563ibus[data_w*1 +:data_w] = c411obus[data_w*4 +:data_w];
assign c411ibus[temp_w*5 +:temp_w] = v1659obus[temp_w*0 +:temp_w];
assign v1659ibus[data_w*0 +:data_w] = c411obus[data_w*5 +:data_w];
assign c412ibus[temp_w*0 +:temp_w] = v259obus[temp_w*2 +:temp_w];
assign v259ibus[data_w*2 +:data_w] = c412obus[data_w*0 +:data_w];
assign c412ibus[temp_w*1 +:temp_w] = v592obus[temp_w*1 +:temp_w];
assign v592ibus[data_w*1 +:data_w] = c412obus[data_w*1 +:data_w];
assign c412ibus[temp_w*2 +:temp_w] = v933obus[temp_w*2 +:temp_w];
assign v933ibus[data_w*2 +:data_w] = c412obus[data_w*2 +:data_w];
assign c412ibus[temp_w*3 +:temp_w] = v964obus[temp_w*0 +:temp_w];
assign v964ibus[data_w*0 +:data_w] = c412obus[data_w*3 +:data_w];
assign c412ibus[temp_w*4 +:temp_w] = v1564obus[temp_w*1 +:temp_w];
assign v1564ibus[data_w*1 +:data_w] = c412obus[data_w*4 +:data_w];
assign c412ibus[temp_w*5 +:temp_w] = v1660obus[temp_w*0 +:temp_w];
assign v1660ibus[data_w*0 +:data_w] = c412obus[data_w*5 +:data_w];
assign c413ibus[temp_w*0 +:temp_w] = v260obus[temp_w*2 +:temp_w];
assign v260ibus[data_w*2 +:data_w] = c413obus[data_w*0 +:data_w];
assign c413ibus[temp_w*1 +:temp_w] = v593obus[temp_w*1 +:temp_w];
assign v593ibus[data_w*1 +:data_w] = c413obus[data_w*1 +:data_w];
assign c413ibus[temp_w*2 +:temp_w] = v934obus[temp_w*2 +:temp_w];
assign v934ibus[data_w*2 +:data_w] = c413obus[data_w*2 +:data_w];
assign c413ibus[temp_w*3 +:temp_w] = v965obus[temp_w*0 +:temp_w];
assign v965ibus[data_w*0 +:data_w] = c413obus[data_w*3 +:data_w];
assign c413ibus[temp_w*4 +:temp_w] = v1565obus[temp_w*1 +:temp_w];
assign v1565ibus[data_w*1 +:data_w] = c413obus[data_w*4 +:data_w];
assign c413ibus[temp_w*5 +:temp_w] = v1661obus[temp_w*0 +:temp_w];
assign v1661ibus[data_w*0 +:data_w] = c413obus[data_w*5 +:data_w];
assign c414ibus[temp_w*0 +:temp_w] = v261obus[temp_w*2 +:temp_w];
assign v261ibus[data_w*2 +:data_w] = c414obus[data_w*0 +:data_w];
assign c414ibus[temp_w*1 +:temp_w] = v594obus[temp_w*1 +:temp_w];
assign v594ibus[data_w*1 +:data_w] = c414obus[data_w*1 +:data_w];
assign c414ibus[temp_w*2 +:temp_w] = v935obus[temp_w*2 +:temp_w];
assign v935ibus[data_w*2 +:data_w] = c414obus[data_w*2 +:data_w];
assign c414ibus[temp_w*3 +:temp_w] = v966obus[temp_w*0 +:temp_w];
assign v966ibus[data_w*0 +:data_w] = c414obus[data_w*3 +:data_w];
assign c414ibus[temp_w*4 +:temp_w] = v1566obus[temp_w*1 +:temp_w];
assign v1566ibus[data_w*1 +:data_w] = c414obus[data_w*4 +:data_w];
assign c414ibus[temp_w*5 +:temp_w] = v1662obus[temp_w*0 +:temp_w];
assign v1662ibus[data_w*0 +:data_w] = c414obus[data_w*5 +:data_w];
assign c415ibus[temp_w*0 +:temp_w] = v262obus[temp_w*2 +:temp_w];
assign v262ibus[data_w*2 +:data_w] = c415obus[data_w*0 +:data_w];
assign c415ibus[temp_w*1 +:temp_w] = v595obus[temp_w*1 +:temp_w];
assign v595ibus[data_w*1 +:data_w] = c415obus[data_w*1 +:data_w];
assign c415ibus[temp_w*2 +:temp_w] = v936obus[temp_w*2 +:temp_w];
assign v936ibus[data_w*2 +:data_w] = c415obus[data_w*2 +:data_w];
assign c415ibus[temp_w*3 +:temp_w] = v967obus[temp_w*0 +:temp_w];
assign v967ibus[data_w*0 +:data_w] = c415obus[data_w*3 +:data_w];
assign c415ibus[temp_w*4 +:temp_w] = v1567obus[temp_w*1 +:temp_w];
assign v1567ibus[data_w*1 +:data_w] = c415obus[data_w*4 +:data_w];
assign c415ibus[temp_w*5 +:temp_w] = v1663obus[temp_w*0 +:temp_w];
assign v1663ibus[data_w*0 +:data_w] = c415obus[data_w*5 +:data_w];
assign c416ibus[temp_w*0 +:temp_w] = v263obus[temp_w*2 +:temp_w];
assign v263ibus[data_w*2 +:data_w] = c416obus[data_w*0 +:data_w];
assign c416ibus[temp_w*1 +:temp_w] = v596obus[temp_w*1 +:temp_w];
assign v596ibus[data_w*1 +:data_w] = c416obus[data_w*1 +:data_w];
assign c416ibus[temp_w*2 +:temp_w] = v937obus[temp_w*2 +:temp_w];
assign v937ibus[data_w*2 +:data_w] = c416obus[data_w*2 +:data_w];
assign c416ibus[temp_w*3 +:temp_w] = v968obus[temp_w*0 +:temp_w];
assign v968ibus[data_w*0 +:data_w] = c416obus[data_w*3 +:data_w];
assign c416ibus[temp_w*4 +:temp_w] = v1568obus[temp_w*1 +:temp_w];
assign v1568ibus[data_w*1 +:data_w] = c416obus[data_w*4 +:data_w];
assign c416ibus[temp_w*5 +:temp_w] = v1664obus[temp_w*0 +:temp_w];
assign v1664ibus[data_w*0 +:data_w] = c416obus[data_w*5 +:data_w];
assign c417ibus[temp_w*0 +:temp_w] = v264obus[temp_w*2 +:temp_w];
assign v264ibus[data_w*2 +:data_w] = c417obus[data_w*0 +:data_w];
assign c417ibus[temp_w*1 +:temp_w] = v597obus[temp_w*1 +:temp_w];
assign v597ibus[data_w*1 +:data_w] = c417obus[data_w*1 +:data_w];
assign c417ibus[temp_w*2 +:temp_w] = v938obus[temp_w*2 +:temp_w];
assign v938ibus[data_w*2 +:data_w] = c417obus[data_w*2 +:data_w];
assign c417ibus[temp_w*3 +:temp_w] = v969obus[temp_w*0 +:temp_w];
assign v969ibus[data_w*0 +:data_w] = c417obus[data_w*3 +:data_w];
assign c417ibus[temp_w*4 +:temp_w] = v1569obus[temp_w*1 +:temp_w];
assign v1569ibus[data_w*1 +:data_w] = c417obus[data_w*4 +:data_w];
assign c417ibus[temp_w*5 +:temp_w] = v1665obus[temp_w*0 +:temp_w];
assign v1665ibus[data_w*0 +:data_w] = c417obus[data_w*5 +:data_w];
assign c418ibus[temp_w*0 +:temp_w] = v265obus[temp_w*2 +:temp_w];
assign v265ibus[data_w*2 +:data_w] = c418obus[data_w*0 +:data_w];
assign c418ibus[temp_w*1 +:temp_w] = v598obus[temp_w*1 +:temp_w];
assign v598ibus[data_w*1 +:data_w] = c418obus[data_w*1 +:data_w];
assign c418ibus[temp_w*2 +:temp_w] = v939obus[temp_w*2 +:temp_w];
assign v939ibus[data_w*2 +:data_w] = c418obus[data_w*2 +:data_w];
assign c418ibus[temp_w*3 +:temp_w] = v970obus[temp_w*0 +:temp_w];
assign v970ibus[data_w*0 +:data_w] = c418obus[data_w*3 +:data_w];
assign c418ibus[temp_w*4 +:temp_w] = v1570obus[temp_w*1 +:temp_w];
assign v1570ibus[data_w*1 +:data_w] = c418obus[data_w*4 +:data_w];
assign c418ibus[temp_w*5 +:temp_w] = v1666obus[temp_w*0 +:temp_w];
assign v1666ibus[data_w*0 +:data_w] = c418obus[data_w*5 +:data_w];
assign c419ibus[temp_w*0 +:temp_w] = v266obus[temp_w*2 +:temp_w];
assign v266ibus[data_w*2 +:data_w] = c419obus[data_w*0 +:data_w];
assign c419ibus[temp_w*1 +:temp_w] = v599obus[temp_w*1 +:temp_w];
assign v599ibus[data_w*1 +:data_w] = c419obus[data_w*1 +:data_w];
assign c419ibus[temp_w*2 +:temp_w] = v940obus[temp_w*2 +:temp_w];
assign v940ibus[data_w*2 +:data_w] = c419obus[data_w*2 +:data_w];
assign c419ibus[temp_w*3 +:temp_w] = v971obus[temp_w*0 +:temp_w];
assign v971ibus[data_w*0 +:data_w] = c419obus[data_w*3 +:data_w];
assign c419ibus[temp_w*4 +:temp_w] = v1571obus[temp_w*1 +:temp_w];
assign v1571ibus[data_w*1 +:data_w] = c419obus[data_w*4 +:data_w];
assign c419ibus[temp_w*5 +:temp_w] = v1667obus[temp_w*0 +:temp_w];
assign v1667ibus[data_w*0 +:data_w] = c419obus[data_w*5 +:data_w];
assign c420ibus[temp_w*0 +:temp_w] = v267obus[temp_w*2 +:temp_w];
assign v267ibus[data_w*2 +:data_w] = c420obus[data_w*0 +:data_w];
assign c420ibus[temp_w*1 +:temp_w] = v600obus[temp_w*1 +:temp_w];
assign v600ibus[data_w*1 +:data_w] = c420obus[data_w*1 +:data_w];
assign c420ibus[temp_w*2 +:temp_w] = v941obus[temp_w*2 +:temp_w];
assign v941ibus[data_w*2 +:data_w] = c420obus[data_w*2 +:data_w];
assign c420ibus[temp_w*3 +:temp_w] = v972obus[temp_w*0 +:temp_w];
assign v972ibus[data_w*0 +:data_w] = c420obus[data_w*3 +:data_w];
assign c420ibus[temp_w*4 +:temp_w] = v1572obus[temp_w*1 +:temp_w];
assign v1572ibus[data_w*1 +:data_w] = c420obus[data_w*4 +:data_w];
assign c420ibus[temp_w*5 +:temp_w] = v1668obus[temp_w*0 +:temp_w];
assign v1668ibus[data_w*0 +:data_w] = c420obus[data_w*5 +:data_w];
assign c421ibus[temp_w*0 +:temp_w] = v268obus[temp_w*2 +:temp_w];
assign v268ibus[data_w*2 +:data_w] = c421obus[data_w*0 +:data_w];
assign c421ibus[temp_w*1 +:temp_w] = v601obus[temp_w*1 +:temp_w];
assign v601ibus[data_w*1 +:data_w] = c421obus[data_w*1 +:data_w];
assign c421ibus[temp_w*2 +:temp_w] = v942obus[temp_w*2 +:temp_w];
assign v942ibus[data_w*2 +:data_w] = c421obus[data_w*2 +:data_w];
assign c421ibus[temp_w*3 +:temp_w] = v973obus[temp_w*0 +:temp_w];
assign v973ibus[data_w*0 +:data_w] = c421obus[data_w*3 +:data_w];
assign c421ibus[temp_w*4 +:temp_w] = v1573obus[temp_w*1 +:temp_w];
assign v1573ibus[data_w*1 +:data_w] = c421obus[data_w*4 +:data_w];
assign c421ibus[temp_w*5 +:temp_w] = v1669obus[temp_w*0 +:temp_w];
assign v1669ibus[data_w*0 +:data_w] = c421obus[data_w*5 +:data_w];
assign c422ibus[temp_w*0 +:temp_w] = v269obus[temp_w*2 +:temp_w];
assign v269ibus[data_w*2 +:data_w] = c422obus[data_w*0 +:data_w];
assign c422ibus[temp_w*1 +:temp_w] = v602obus[temp_w*1 +:temp_w];
assign v602ibus[data_w*1 +:data_w] = c422obus[data_w*1 +:data_w];
assign c422ibus[temp_w*2 +:temp_w] = v943obus[temp_w*2 +:temp_w];
assign v943ibus[data_w*2 +:data_w] = c422obus[data_w*2 +:data_w];
assign c422ibus[temp_w*3 +:temp_w] = v974obus[temp_w*0 +:temp_w];
assign v974ibus[data_w*0 +:data_w] = c422obus[data_w*3 +:data_w];
assign c422ibus[temp_w*4 +:temp_w] = v1574obus[temp_w*1 +:temp_w];
assign v1574ibus[data_w*1 +:data_w] = c422obus[data_w*4 +:data_w];
assign c422ibus[temp_w*5 +:temp_w] = v1670obus[temp_w*0 +:temp_w];
assign v1670ibus[data_w*0 +:data_w] = c422obus[data_w*5 +:data_w];
assign c423ibus[temp_w*0 +:temp_w] = v270obus[temp_w*2 +:temp_w];
assign v270ibus[data_w*2 +:data_w] = c423obus[data_w*0 +:data_w];
assign c423ibus[temp_w*1 +:temp_w] = v603obus[temp_w*1 +:temp_w];
assign v603ibus[data_w*1 +:data_w] = c423obus[data_w*1 +:data_w];
assign c423ibus[temp_w*2 +:temp_w] = v944obus[temp_w*2 +:temp_w];
assign v944ibus[data_w*2 +:data_w] = c423obus[data_w*2 +:data_w];
assign c423ibus[temp_w*3 +:temp_w] = v975obus[temp_w*0 +:temp_w];
assign v975ibus[data_w*0 +:data_w] = c423obus[data_w*3 +:data_w];
assign c423ibus[temp_w*4 +:temp_w] = v1575obus[temp_w*1 +:temp_w];
assign v1575ibus[data_w*1 +:data_w] = c423obus[data_w*4 +:data_w];
assign c423ibus[temp_w*5 +:temp_w] = v1671obus[temp_w*0 +:temp_w];
assign v1671ibus[data_w*0 +:data_w] = c423obus[data_w*5 +:data_w];
assign c424ibus[temp_w*0 +:temp_w] = v271obus[temp_w*2 +:temp_w];
assign v271ibus[data_w*2 +:data_w] = c424obus[data_w*0 +:data_w];
assign c424ibus[temp_w*1 +:temp_w] = v604obus[temp_w*1 +:temp_w];
assign v604ibus[data_w*1 +:data_w] = c424obus[data_w*1 +:data_w];
assign c424ibus[temp_w*2 +:temp_w] = v945obus[temp_w*2 +:temp_w];
assign v945ibus[data_w*2 +:data_w] = c424obus[data_w*2 +:data_w];
assign c424ibus[temp_w*3 +:temp_w] = v976obus[temp_w*0 +:temp_w];
assign v976ibus[data_w*0 +:data_w] = c424obus[data_w*3 +:data_w];
assign c424ibus[temp_w*4 +:temp_w] = v1576obus[temp_w*1 +:temp_w];
assign v1576ibus[data_w*1 +:data_w] = c424obus[data_w*4 +:data_w];
assign c424ibus[temp_w*5 +:temp_w] = v1672obus[temp_w*0 +:temp_w];
assign v1672ibus[data_w*0 +:data_w] = c424obus[data_w*5 +:data_w];
assign c425ibus[temp_w*0 +:temp_w] = v272obus[temp_w*2 +:temp_w];
assign v272ibus[data_w*2 +:data_w] = c425obus[data_w*0 +:data_w];
assign c425ibus[temp_w*1 +:temp_w] = v605obus[temp_w*1 +:temp_w];
assign v605ibus[data_w*1 +:data_w] = c425obus[data_w*1 +:data_w];
assign c425ibus[temp_w*2 +:temp_w] = v946obus[temp_w*2 +:temp_w];
assign v946ibus[data_w*2 +:data_w] = c425obus[data_w*2 +:data_w];
assign c425ibus[temp_w*3 +:temp_w] = v977obus[temp_w*0 +:temp_w];
assign v977ibus[data_w*0 +:data_w] = c425obus[data_w*3 +:data_w];
assign c425ibus[temp_w*4 +:temp_w] = v1577obus[temp_w*1 +:temp_w];
assign v1577ibus[data_w*1 +:data_w] = c425obus[data_w*4 +:data_w];
assign c425ibus[temp_w*5 +:temp_w] = v1673obus[temp_w*0 +:temp_w];
assign v1673ibus[data_w*0 +:data_w] = c425obus[data_w*5 +:data_w];
assign c426ibus[temp_w*0 +:temp_w] = v273obus[temp_w*2 +:temp_w];
assign v273ibus[data_w*2 +:data_w] = c426obus[data_w*0 +:data_w];
assign c426ibus[temp_w*1 +:temp_w] = v606obus[temp_w*1 +:temp_w];
assign v606ibus[data_w*1 +:data_w] = c426obus[data_w*1 +:data_w];
assign c426ibus[temp_w*2 +:temp_w] = v947obus[temp_w*2 +:temp_w];
assign v947ibus[data_w*2 +:data_w] = c426obus[data_w*2 +:data_w];
assign c426ibus[temp_w*3 +:temp_w] = v978obus[temp_w*0 +:temp_w];
assign v978ibus[data_w*0 +:data_w] = c426obus[data_w*3 +:data_w];
assign c426ibus[temp_w*4 +:temp_w] = v1578obus[temp_w*1 +:temp_w];
assign v1578ibus[data_w*1 +:data_w] = c426obus[data_w*4 +:data_w];
assign c426ibus[temp_w*5 +:temp_w] = v1674obus[temp_w*0 +:temp_w];
assign v1674ibus[data_w*0 +:data_w] = c426obus[data_w*5 +:data_w];
assign c427ibus[temp_w*0 +:temp_w] = v274obus[temp_w*2 +:temp_w];
assign v274ibus[data_w*2 +:data_w] = c427obus[data_w*0 +:data_w];
assign c427ibus[temp_w*1 +:temp_w] = v607obus[temp_w*1 +:temp_w];
assign v607ibus[data_w*1 +:data_w] = c427obus[data_w*1 +:data_w];
assign c427ibus[temp_w*2 +:temp_w] = v948obus[temp_w*2 +:temp_w];
assign v948ibus[data_w*2 +:data_w] = c427obus[data_w*2 +:data_w];
assign c427ibus[temp_w*3 +:temp_w] = v979obus[temp_w*0 +:temp_w];
assign v979ibus[data_w*0 +:data_w] = c427obus[data_w*3 +:data_w];
assign c427ibus[temp_w*4 +:temp_w] = v1579obus[temp_w*1 +:temp_w];
assign v1579ibus[data_w*1 +:data_w] = c427obus[data_w*4 +:data_w];
assign c427ibus[temp_w*5 +:temp_w] = v1675obus[temp_w*0 +:temp_w];
assign v1675ibus[data_w*0 +:data_w] = c427obus[data_w*5 +:data_w];
assign c428ibus[temp_w*0 +:temp_w] = v275obus[temp_w*2 +:temp_w];
assign v275ibus[data_w*2 +:data_w] = c428obus[data_w*0 +:data_w];
assign c428ibus[temp_w*1 +:temp_w] = v608obus[temp_w*1 +:temp_w];
assign v608ibus[data_w*1 +:data_w] = c428obus[data_w*1 +:data_w];
assign c428ibus[temp_w*2 +:temp_w] = v949obus[temp_w*2 +:temp_w];
assign v949ibus[data_w*2 +:data_w] = c428obus[data_w*2 +:data_w];
assign c428ibus[temp_w*3 +:temp_w] = v980obus[temp_w*0 +:temp_w];
assign v980ibus[data_w*0 +:data_w] = c428obus[data_w*3 +:data_w];
assign c428ibus[temp_w*4 +:temp_w] = v1580obus[temp_w*1 +:temp_w];
assign v1580ibus[data_w*1 +:data_w] = c428obus[data_w*4 +:data_w];
assign c428ibus[temp_w*5 +:temp_w] = v1676obus[temp_w*0 +:temp_w];
assign v1676ibus[data_w*0 +:data_w] = c428obus[data_w*5 +:data_w];
assign c429ibus[temp_w*0 +:temp_w] = v276obus[temp_w*2 +:temp_w];
assign v276ibus[data_w*2 +:data_w] = c429obus[data_w*0 +:data_w];
assign c429ibus[temp_w*1 +:temp_w] = v609obus[temp_w*1 +:temp_w];
assign v609ibus[data_w*1 +:data_w] = c429obus[data_w*1 +:data_w];
assign c429ibus[temp_w*2 +:temp_w] = v950obus[temp_w*2 +:temp_w];
assign v950ibus[data_w*2 +:data_w] = c429obus[data_w*2 +:data_w];
assign c429ibus[temp_w*3 +:temp_w] = v981obus[temp_w*0 +:temp_w];
assign v981ibus[data_w*0 +:data_w] = c429obus[data_w*3 +:data_w];
assign c429ibus[temp_w*4 +:temp_w] = v1581obus[temp_w*1 +:temp_w];
assign v1581ibus[data_w*1 +:data_w] = c429obus[data_w*4 +:data_w];
assign c429ibus[temp_w*5 +:temp_w] = v1677obus[temp_w*0 +:temp_w];
assign v1677ibus[data_w*0 +:data_w] = c429obus[data_w*5 +:data_w];
assign c430ibus[temp_w*0 +:temp_w] = v277obus[temp_w*2 +:temp_w];
assign v277ibus[data_w*2 +:data_w] = c430obus[data_w*0 +:data_w];
assign c430ibus[temp_w*1 +:temp_w] = v610obus[temp_w*1 +:temp_w];
assign v610ibus[data_w*1 +:data_w] = c430obus[data_w*1 +:data_w];
assign c430ibus[temp_w*2 +:temp_w] = v951obus[temp_w*2 +:temp_w];
assign v951ibus[data_w*2 +:data_w] = c430obus[data_w*2 +:data_w];
assign c430ibus[temp_w*3 +:temp_w] = v982obus[temp_w*0 +:temp_w];
assign v982ibus[data_w*0 +:data_w] = c430obus[data_w*3 +:data_w];
assign c430ibus[temp_w*4 +:temp_w] = v1582obus[temp_w*1 +:temp_w];
assign v1582ibus[data_w*1 +:data_w] = c430obus[data_w*4 +:data_w];
assign c430ibus[temp_w*5 +:temp_w] = v1678obus[temp_w*0 +:temp_w];
assign v1678ibus[data_w*0 +:data_w] = c430obus[data_w*5 +:data_w];
assign c431ibus[temp_w*0 +:temp_w] = v278obus[temp_w*2 +:temp_w];
assign v278ibus[data_w*2 +:data_w] = c431obus[data_w*0 +:data_w];
assign c431ibus[temp_w*1 +:temp_w] = v611obus[temp_w*1 +:temp_w];
assign v611ibus[data_w*1 +:data_w] = c431obus[data_w*1 +:data_w];
assign c431ibus[temp_w*2 +:temp_w] = v952obus[temp_w*2 +:temp_w];
assign v952ibus[data_w*2 +:data_w] = c431obus[data_w*2 +:data_w];
assign c431ibus[temp_w*3 +:temp_w] = v983obus[temp_w*0 +:temp_w];
assign v983ibus[data_w*0 +:data_w] = c431obus[data_w*3 +:data_w];
assign c431ibus[temp_w*4 +:temp_w] = v1583obus[temp_w*1 +:temp_w];
assign v1583ibus[data_w*1 +:data_w] = c431obus[data_w*4 +:data_w];
assign c431ibus[temp_w*5 +:temp_w] = v1679obus[temp_w*0 +:temp_w];
assign v1679ibus[data_w*0 +:data_w] = c431obus[data_w*5 +:data_w];
assign c432ibus[temp_w*0 +:temp_w] = v279obus[temp_w*2 +:temp_w];
assign v279ibus[data_w*2 +:data_w] = c432obus[data_w*0 +:data_w];
assign c432ibus[temp_w*1 +:temp_w] = v612obus[temp_w*1 +:temp_w];
assign v612ibus[data_w*1 +:data_w] = c432obus[data_w*1 +:data_w];
assign c432ibus[temp_w*2 +:temp_w] = v953obus[temp_w*2 +:temp_w];
assign v953ibus[data_w*2 +:data_w] = c432obus[data_w*2 +:data_w];
assign c432ibus[temp_w*3 +:temp_w] = v984obus[temp_w*0 +:temp_w];
assign v984ibus[data_w*0 +:data_w] = c432obus[data_w*3 +:data_w];
assign c432ibus[temp_w*4 +:temp_w] = v1584obus[temp_w*1 +:temp_w];
assign v1584ibus[data_w*1 +:data_w] = c432obus[data_w*4 +:data_w];
assign c432ibus[temp_w*5 +:temp_w] = v1680obus[temp_w*0 +:temp_w];
assign v1680ibus[data_w*0 +:data_w] = c432obus[data_w*5 +:data_w];
assign c433ibus[temp_w*0 +:temp_w] = v280obus[temp_w*2 +:temp_w];
assign v280ibus[data_w*2 +:data_w] = c433obus[data_w*0 +:data_w];
assign c433ibus[temp_w*1 +:temp_w] = v613obus[temp_w*1 +:temp_w];
assign v613ibus[data_w*1 +:data_w] = c433obus[data_w*1 +:data_w];
assign c433ibus[temp_w*2 +:temp_w] = v954obus[temp_w*2 +:temp_w];
assign v954ibus[data_w*2 +:data_w] = c433obus[data_w*2 +:data_w];
assign c433ibus[temp_w*3 +:temp_w] = v985obus[temp_w*0 +:temp_w];
assign v985ibus[data_w*0 +:data_w] = c433obus[data_w*3 +:data_w];
assign c433ibus[temp_w*4 +:temp_w] = v1585obus[temp_w*1 +:temp_w];
assign v1585ibus[data_w*1 +:data_w] = c433obus[data_w*4 +:data_w];
assign c433ibus[temp_w*5 +:temp_w] = v1681obus[temp_w*0 +:temp_w];
assign v1681ibus[data_w*0 +:data_w] = c433obus[data_w*5 +:data_w];
assign c434ibus[temp_w*0 +:temp_w] = v281obus[temp_w*2 +:temp_w];
assign v281ibus[data_w*2 +:data_w] = c434obus[data_w*0 +:data_w];
assign c434ibus[temp_w*1 +:temp_w] = v614obus[temp_w*1 +:temp_w];
assign v614ibus[data_w*1 +:data_w] = c434obus[data_w*1 +:data_w];
assign c434ibus[temp_w*2 +:temp_w] = v955obus[temp_w*2 +:temp_w];
assign v955ibus[data_w*2 +:data_w] = c434obus[data_w*2 +:data_w];
assign c434ibus[temp_w*3 +:temp_w] = v986obus[temp_w*0 +:temp_w];
assign v986ibus[data_w*0 +:data_w] = c434obus[data_w*3 +:data_w];
assign c434ibus[temp_w*4 +:temp_w] = v1586obus[temp_w*1 +:temp_w];
assign v1586ibus[data_w*1 +:data_w] = c434obus[data_w*4 +:data_w];
assign c434ibus[temp_w*5 +:temp_w] = v1682obus[temp_w*0 +:temp_w];
assign v1682ibus[data_w*0 +:data_w] = c434obus[data_w*5 +:data_w];
assign c435ibus[temp_w*0 +:temp_w] = v282obus[temp_w*2 +:temp_w];
assign v282ibus[data_w*2 +:data_w] = c435obus[data_w*0 +:data_w];
assign c435ibus[temp_w*1 +:temp_w] = v615obus[temp_w*1 +:temp_w];
assign v615ibus[data_w*1 +:data_w] = c435obus[data_w*1 +:data_w];
assign c435ibus[temp_w*2 +:temp_w] = v956obus[temp_w*2 +:temp_w];
assign v956ibus[data_w*2 +:data_w] = c435obus[data_w*2 +:data_w];
assign c435ibus[temp_w*3 +:temp_w] = v987obus[temp_w*0 +:temp_w];
assign v987ibus[data_w*0 +:data_w] = c435obus[data_w*3 +:data_w];
assign c435ibus[temp_w*4 +:temp_w] = v1587obus[temp_w*1 +:temp_w];
assign v1587ibus[data_w*1 +:data_w] = c435obus[data_w*4 +:data_w];
assign c435ibus[temp_w*5 +:temp_w] = v1683obus[temp_w*0 +:temp_w];
assign v1683ibus[data_w*0 +:data_w] = c435obus[data_w*5 +:data_w];
assign c436ibus[temp_w*0 +:temp_w] = v283obus[temp_w*2 +:temp_w];
assign v283ibus[data_w*2 +:data_w] = c436obus[data_w*0 +:data_w];
assign c436ibus[temp_w*1 +:temp_w] = v616obus[temp_w*1 +:temp_w];
assign v616ibus[data_w*1 +:data_w] = c436obus[data_w*1 +:data_w];
assign c436ibus[temp_w*2 +:temp_w] = v957obus[temp_w*2 +:temp_w];
assign v957ibus[data_w*2 +:data_w] = c436obus[data_w*2 +:data_w];
assign c436ibus[temp_w*3 +:temp_w] = v988obus[temp_w*0 +:temp_w];
assign v988ibus[data_w*0 +:data_w] = c436obus[data_w*3 +:data_w];
assign c436ibus[temp_w*4 +:temp_w] = v1588obus[temp_w*1 +:temp_w];
assign v1588ibus[data_w*1 +:data_w] = c436obus[data_w*4 +:data_w];
assign c436ibus[temp_w*5 +:temp_w] = v1684obus[temp_w*0 +:temp_w];
assign v1684ibus[data_w*0 +:data_w] = c436obus[data_w*5 +:data_w];
assign c437ibus[temp_w*0 +:temp_w] = v284obus[temp_w*2 +:temp_w];
assign v284ibus[data_w*2 +:data_w] = c437obus[data_w*0 +:data_w];
assign c437ibus[temp_w*1 +:temp_w] = v617obus[temp_w*1 +:temp_w];
assign v617ibus[data_w*1 +:data_w] = c437obus[data_w*1 +:data_w];
assign c437ibus[temp_w*2 +:temp_w] = v958obus[temp_w*2 +:temp_w];
assign v958ibus[data_w*2 +:data_w] = c437obus[data_w*2 +:data_w];
assign c437ibus[temp_w*3 +:temp_w] = v989obus[temp_w*0 +:temp_w];
assign v989ibus[data_w*0 +:data_w] = c437obus[data_w*3 +:data_w];
assign c437ibus[temp_w*4 +:temp_w] = v1589obus[temp_w*1 +:temp_w];
assign v1589ibus[data_w*1 +:data_w] = c437obus[data_w*4 +:data_w];
assign c437ibus[temp_w*5 +:temp_w] = v1685obus[temp_w*0 +:temp_w];
assign v1685ibus[data_w*0 +:data_w] = c437obus[data_w*5 +:data_w];
assign c438ibus[temp_w*0 +:temp_w] = v285obus[temp_w*2 +:temp_w];
assign v285ibus[data_w*2 +:data_w] = c438obus[data_w*0 +:data_w];
assign c438ibus[temp_w*1 +:temp_w] = v618obus[temp_w*1 +:temp_w];
assign v618ibus[data_w*1 +:data_w] = c438obus[data_w*1 +:data_w];
assign c438ibus[temp_w*2 +:temp_w] = v959obus[temp_w*2 +:temp_w];
assign v959ibus[data_w*2 +:data_w] = c438obus[data_w*2 +:data_w];
assign c438ibus[temp_w*3 +:temp_w] = v990obus[temp_w*0 +:temp_w];
assign v990ibus[data_w*0 +:data_w] = c438obus[data_w*3 +:data_w];
assign c438ibus[temp_w*4 +:temp_w] = v1590obus[temp_w*1 +:temp_w];
assign v1590ibus[data_w*1 +:data_w] = c438obus[data_w*4 +:data_w];
assign c438ibus[temp_w*5 +:temp_w] = v1686obus[temp_w*0 +:temp_w];
assign v1686ibus[data_w*0 +:data_w] = c438obus[data_w*5 +:data_w];
assign c439ibus[temp_w*0 +:temp_w] = v286obus[temp_w*2 +:temp_w];
assign v286ibus[data_w*2 +:data_w] = c439obus[data_w*0 +:data_w];
assign c439ibus[temp_w*1 +:temp_w] = v619obus[temp_w*1 +:temp_w];
assign v619ibus[data_w*1 +:data_w] = c439obus[data_w*1 +:data_w];
assign c439ibus[temp_w*2 +:temp_w] = v864obus[temp_w*2 +:temp_w];
assign v864ibus[data_w*2 +:data_w] = c439obus[data_w*2 +:data_w];
assign c439ibus[temp_w*3 +:temp_w] = v991obus[temp_w*0 +:temp_w];
assign v991ibus[data_w*0 +:data_w] = c439obus[data_w*3 +:data_w];
assign c439ibus[temp_w*4 +:temp_w] = v1591obus[temp_w*1 +:temp_w];
assign v1591ibus[data_w*1 +:data_w] = c439obus[data_w*4 +:data_w];
assign c439ibus[temp_w*5 +:temp_w] = v1687obus[temp_w*0 +:temp_w];
assign v1687ibus[data_w*0 +:data_w] = c439obus[data_w*5 +:data_w];
assign c440ibus[temp_w*0 +:temp_w] = v287obus[temp_w*2 +:temp_w];
assign v287ibus[data_w*2 +:data_w] = c440obus[data_w*0 +:data_w];
assign c440ibus[temp_w*1 +:temp_w] = v620obus[temp_w*1 +:temp_w];
assign v620ibus[data_w*1 +:data_w] = c440obus[data_w*1 +:data_w];
assign c440ibus[temp_w*2 +:temp_w] = v865obus[temp_w*2 +:temp_w];
assign v865ibus[data_w*2 +:data_w] = c440obus[data_w*2 +:data_w];
assign c440ibus[temp_w*3 +:temp_w] = v992obus[temp_w*0 +:temp_w];
assign v992ibus[data_w*0 +:data_w] = c440obus[data_w*3 +:data_w];
assign c440ibus[temp_w*4 +:temp_w] = v1592obus[temp_w*1 +:temp_w];
assign v1592ibus[data_w*1 +:data_w] = c440obus[data_w*4 +:data_w];
assign c440ibus[temp_w*5 +:temp_w] = v1688obus[temp_w*0 +:temp_w];
assign v1688ibus[data_w*0 +:data_w] = c440obus[data_w*5 +:data_w];
assign c441ibus[temp_w*0 +:temp_w] = v192obus[temp_w*2 +:temp_w];
assign v192ibus[data_w*2 +:data_w] = c441obus[data_w*0 +:data_w];
assign c441ibus[temp_w*1 +:temp_w] = v621obus[temp_w*1 +:temp_w];
assign v621ibus[data_w*1 +:data_w] = c441obus[data_w*1 +:data_w];
assign c441ibus[temp_w*2 +:temp_w] = v866obus[temp_w*2 +:temp_w];
assign v866ibus[data_w*2 +:data_w] = c441obus[data_w*2 +:data_w];
assign c441ibus[temp_w*3 +:temp_w] = v993obus[temp_w*0 +:temp_w];
assign v993ibus[data_w*0 +:data_w] = c441obus[data_w*3 +:data_w];
assign c441ibus[temp_w*4 +:temp_w] = v1593obus[temp_w*1 +:temp_w];
assign v1593ibus[data_w*1 +:data_w] = c441obus[data_w*4 +:data_w];
assign c441ibus[temp_w*5 +:temp_w] = v1689obus[temp_w*0 +:temp_w];
assign v1689ibus[data_w*0 +:data_w] = c441obus[data_w*5 +:data_w];
assign c442ibus[temp_w*0 +:temp_w] = v193obus[temp_w*2 +:temp_w];
assign v193ibus[data_w*2 +:data_w] = c442obus[data_w*0 +:data_w];
assign c442ibus[temp_w*1 +:temp_w] = v622obus[temp_w*1 +:temp_w];
assign v622ibus[data_w*1 +:data_w] = c442obus[data_w*1 +:data_w];
assign c442ibus[temp_w*2 +:temp_w] = v867obus[temp_w*2 +:temp_w];
assign v867ibus[data_w*2 +:data_w] = c442obus[data_w*2 +:data_w];
assign c442ibus[temp_w*3 +:temp_w] = v994obus[temp_w*0 +:temp_w];
assign v994ibus[data_w*0 +:data_w] = c442obus[data_w*3 +:data_w];
assign c442ibus[temp_w*4 +:temp_w] = v1594obus[temp_w*1 +:temp_w];
assign v1594ibus[data_w*1 +:data_w] = c442obus[data_w*4 +:data_w];
assign c442ibus[temp_w*5 +:temp_w] = v1690obus[temp_w*0 +:temp_w];
assign v1690ibus[data_w*0 +:data_w] = c442obus[data_w*5 +:data_w];
assign c443ibus[temp_w*0 +:temp_w] = v194obus[temp_w*2 +:temp_w];
assign v194ibus[data_w*2 +:data_w] = c443obus[data_w*0 +:data_w];
assign c443ibus[temp_w*1 +:temp_w] = v623obus[temp_w*1 +:temp_w];
assign v623ibus[data_w*1 +:data_w] = c443obus[data_w*1 +:data_w];
assign c443ibus[temp_w*2 +:temp_w] = v868obus[temp_w*2 +:temp_w];
assign v868ibus[data_w*2 +:data_w] = c443obus[data_w*2 +:data_w];
assign c443ibus[temp_w*3 +:temp_w] = v995obus[temp_w*0 +:temp_w];
assign v995ibus[data_w*0 +:data_w] = c443obus[data_w*3 +:data_w];
assign c443ibus[temp_w*4 +:temp_w] = v1595obus[temp_w*1 +:temp_w];
assign v1595ibus[data_w*1 +:data_w] = c443obus[data_w*4 +:data_w];
assign c443ibus[temp_w*5 +:temp_w] = v1691obus[temp_w*0 +:temp_w];
assign v1691ibus[data_w*0 +:data_w] = c443obus[data_w*5 +:data_w];
assign c444ibus[temp_w*0 +:temp_w] = v195obus[temp_w*2 +:temp_w];
assign v195ibus[data_w*2 +:data_w] = c444obus[data_w*0 +:data_w];
assign c444ibus[temp_w*1 +:temp_w] = v624obus[temp_w*1 +:temp_w];
assign v624ibus[data_w*1 +:data_w] = c444obus[data_w*1 +:data_w];
assign c444ibus[temp_w*2 +:temp_w] = v869obus[temp_w*2 +:temp_w];
assign v869ibus[data_w*2 +:data_w] = c444obus[data_w*2 +:data_w];
assign c444ibus[temp_w*3 +:temp_w] = v996obus[temp_w*0 +:temp_w];
assign v996ibus[data_w*0 +:data_w] = c444obus[data_w*3 +:data_w];
assign c444ibus[temp_w*4 +:temp_w] = v1596obus[temp_w*1 +:temp_w];
assign v1596ibus[data_w*1 +:data_w] = c444obus[data_w*4 +:data_w];
assign c444ibus[temp_w*5 +:temp_w] = v1692obus[temp_w*0 +:temp_w];
assign v1692ibus[data_w*0 +:data_w] = c444obus[data_w*5 +:data_w];
assign c445ibus[temp_w*0 +:temp_w] = v196obus[temp_w*2 +:temp_w];
assign v196ibus[data_w*2 +:data_w] = c445obus[data_w*0 +:data_w];
assign c445ibus[temp_w*1 +:temp_w] = v625obus[temp_w*1 +:temp_w];
assign v625ibus[data_w*1 +:data_w] = c445obus[data_w*1 +:data_w];
assign c445ibus[temp_w*2 +:temp_w] = v870obus[temp_w*2 +:temp_w];
assign v870ibus[data_w*2 +:data_w] = c445obus[data_w*2 +:data_w];
assign c445ibus[temp_w*3 +:temp_w] = v997obus[temp_w*0 +:temp_w];
assign v997ibus[data_w*0 +:data_w] = c445obus[data_w*3 +:data_w];
assign c445ibus[temp_w*4 +:temp_w] = v1597obus[temp_w*1 +:temp_w];
assign v1597ibus[data_w*1 +:data_w] = c445obus[data_w*4 +:data_w];
assign c445ibus[temp_w*5 +:temp_w] = v1693obus[temp_w*0 +:temp_w];
assign v1693ibus[data_w*0 +:data_w] = c445obus[data_w*5 +:data_w];
assign c446ibus[temp_w*0 +:temp_w] = v197obus[temp_w*2 +:temp_w];
assign v197ibus[data_w*2 +:data_w] = c446obus[data_w*0 +:data_w];
assign c446ibus[temp_w*1 +:temp_w] = v626obus[temp_w*1 +:temp_w];
assign v626ibus[data_w*1 +:data_w] = c446obus[data_w*1 +:data_w];
assign c446ibus[temp_w*2 +:temp_w] = v871obus[temp_w*2 +:temp_w];
assign v871ibus[data_w*2 +:data_w] = c446obus[data_w*2 +:data_w];
assign c446ibus[temp_w*3 +:temp_w] = v998obus[temp_w*0 +:temp_w];
assign v998ibus[data_w*0 +:data_w] = c446obus[data_w*3 +:data_w];
assign c446ibus[temp_w*4 +:temp_w] = v1598obus[temp_w*1 +:temp_w];
assign v1598ibus[data_w*1 +:data_w] = c446obus[data_w*4 +:data_w];
assign c446ibus[temp_w*5 +:temp_w] = v1694obus[temp_w*0 +:temp_w];
assign v1694ibus[data_w*0 +:data_w] = c446obus[data_w*5 +:data_w];
assign c447ibus[temp_w*0 +:temp_w] = v198obus[temp_w*2 +:temp_w];
assign v198ibus[data_w*2 +:data_w] = c447obus[data_w*0 +:data_w];
assign c447ibus[temp_w*1 +:temp_w] = v627obus[temp_w*1 +:temp_w];
assign v627ibus[data_w*1 +:data_w] = c447obus[data_w*1 +:data_w];
assign c447ibus[temp_w*2 +:temp_w] = v872obus[temp_w*2 +:temp_w];
assign v872ibus[data_w*2 +:data_w] = c447obus[data_w*2 +:data_w];
assign c447ibus[temp_w*3 +:temp_w] = v999obus[temp_w*0 +:temp_w];
assign v999ibus[data_w*0 +:data_w] = c447obus[data_w*3 +:data_w];
assign c447ibus[temp_w*4 +:temp_w] = v1599obus[temp_w*1 +:temp_w];
assign v1599ibus[data_w*1 +:data_w] = c447obus[data_w*4 +:data_w];
assign c447ibus[temp_w*5 +:temp_w] = v1695obus[temp_w*0 +:temp_w];
assign v1695ibus[data_w*0 +:data_w] = c447obus[data_w*5 +:data_w];
assign c448ibus[temp_w*0 +:temp_w] = v199obus[temp_w*2 +:temp_w];
assign v199ibus[data_w*2 +:data_w] = c448obus[data_w*0 +:data_w];
assign c448ibus[temp_w*1 +:temp_w] = v628obus[temp_w*1 +:temp_w];
assign v628ibus[data_w*1 +:data_w] = c448obus[data_w*1 +:data_w];
assign c448ibus[temp_w*2 +:temp_w] = v873obus[temp_w*2 +:temp_w];
assign v873ibus[data_w*2 +:data_w] = c448obus[data_w*2 +:data_w];
assign c448ibus[temp_w*3 +:temp_w] = v1000obus[temp_w*0 +:temp_w];
assign v1000ibus[data_w*0 +:data_w] = c448obus[data_w*3 +:data_w];
assign c448ibus[temp_w*4 +:temp_w] = v1600obus[temp_w*1 +:temp_w];
assign v1600ibus[data_w*1 +:data_w] = c448obus[data_w*4 +:data_w];
assign c448ibus[temp_w*5 +:temp_w] = v1696obus[temp_w*0 +:temp_w];
assign v1696ibus[data_w*0 +:data_w] = c448obus[data_w*5 +:data_w];
assign c449ibus[temp_w*0 +:temp_w] = v200obus[temp_w*2 +:temp_w];
assign v200ibus[data_w*2 +:data_w] = c449obus[data_w*0 +:data_w];
assign c449ibus[temp_w*1 +:temp_w] = v629obus[temp_w*1 +:temp_w];
assign v629ibus[data_w*1 +:data_w] = c449obus[data_w*1 +:data_w];
assign c449ibus[temp_w*2 +:temp_w] = v874obus[temp_w*2 +:temp_w];
assign v874ibus[data_w*2 +:data_w] = c449obus[data_w*2 +:data_w];
assign c449ibus[temp_w*3 +:temp_w] = v1001obus[temp_w*0 +:temp_w];
assign v1001ibus[data_w*0 +:data_w] = c449obus[data_w*3 +:data_w];
assign c449ibus[temp_w*4 +:temp_w] = v1601obus[temp_w*1 +:temp_w];
assign v1601ibus[data_w*1 +:data_w] = c449obus[data_w*4 +:data_w];
assign c449ibus[temp_w*5 +:temp_w] = v1697obus[temp_w*0 +:temp_w];
assign v1697ibus[data_w*0 +:data_w] = c449obus[data_w*5 +:data_w];
assign c450ibus[temp_w*0 +:temp_w] = v201obus[temp_w*2 +:temp_w];
assign v201ibus[data_w*2 +:data_w] = c450obus[data_w*0 +:data_w];
assign c450ibus[temp_w*1 +:temp_w] = v630obus[temp_w*1 +:temp_w];
assign v630ibus[data_w*1 +:data_w] = c450obus[data_w*1 +:data_w];
assign c450ibus[temp_w*2 +:temp_w] = v875obus[temp_w*2 +:temp_w];
assign v875ibus[data_w*2 +:data_w] = c450obus[data_w*2 +:data_w];
assign c450ibus[temp_w*3 +:temp_w] = v1002obus[temp_w*0 +:temp_w];
assign v1002ibus[data_w*0 +:data_w] = c450obus[data_w*3 +:data_w];
assign c450ibus[temp_w*4 +:temp_w] = v1602obus[temp_w*1 +:temp_w];
assign v1602ibus[data_w*1 +:data_w] = c450obus[data_w*4 +:data_w];
assign c450ibus[temp_w*5 +:temp_w] = v1698obus[temp_w*0 +:temp_w];
assign v1698ibus[data_w*0 +:data_w] = c450obus[data_w*5 +:data_w];
assign c451ibus[temp_w*0 +:temp_w] = v202obus[temp_w*2 +:temp_w];
assign v202ibus[data_w*2 +:data_w] = c451obus[data_w*0 +:data_w];
assign c451ibus[temp_w*1 +:temp_w] = v631obus[temp_w*1 +:temp_w];
assign v631ibus[data_w*1 +:data_w] = c451obus[data_w*1 +:data_w];
assign c451ibus[temp_w*2 +:temp_w] = v876obus[temp_w*2 +:temp_w];
assign v876ibus[data_w*2 +:data_w] = c451obus[data_w*2 +:data_w];
assign c451ibus[temp_w*3 +:temp_w] = v1003obus[temp_w*0 +:temp_w];
assign v1003ibus[data_w*0 +:data_w] = c451obus[data_w*3 +:data_w];
assign c451ibus[temp_w*4 +:temp_w] = v1603obus[temp_w*1 +:temp_w];
assign v1603ibus[data_w*1 +:data_w] = c451obus[data_w*4 +:data_w];
assign c451ibus[temp_w*5 +:temp_w] = v1699obus[temp_w*0 +:temp_w];
assign v1699ibus[data_w*0 +:data_w] = c451obus[data_w*5 +:data_w];
assign c452ibus[temp_w*0 +:temp_w] = v203obus[temp_w*2 +:temp_w];
assign v203ibus[data_w*2 +:data_w] = c452obus[data_w*0 +:data_w];
assign c452ibus[temp_w*1 +:temp_w] = v632obus[temp_w*1 +:temp_w];
assign v632ibus[data_w*1 +:data_w] = c452obus[data_w*1 +:data_w];
assign c452ibus[temp_w*2 +:temp_w] = v877obus[temp_w*2 +:temp_w];
assign v877ibus[data_w*2 +:data_w] = c452obus[data_w*2 +:data_w];
assign c452ibus[temp_w*3 +:temp_w] = v1004obus[temp_w*0 +:temp_w];
assign v1004ibus[data_w*0 +:data_w] = c452obus[data_w*3 +:data_w];
assign c452ibus[temp_w*4 +:temp_w] = v1604obus[temp_w*1 +:temp_w];
assign v1604ibus[data_w*1 +:data_w] = c452obus[data_w*4 +:data_w];
assign c452ibus[temp_w*5 +:temp_w] = v1700obus[temp_w*0 +:temp_w];
assign v1700ibus[data_w*0 +:data_w] = c452obus[data_w*5 +:data_w];
assign c453ibus[temp_w*0 +:temp_w] = v204obus[temp_w*2 +:temp_w];
assign v204ibus[data_w*2 +:data_w] = c453obus[data_w*0 +:data_w];
assign c453ibus[temp_w*1 +:temp_w] = v633obus[temp_w*1 +:temp_w];
assign v633ibus[data_w*1 +:data_w] = c453obus[data_w*1 +:data_w];
assign c453ibus[temp_w*2 +:temp_w] = v878obus[temp_w*2 +:temp_w];
assign v878ibus[data_w*2 +:data_w] = c453obus[data_w*2 +:data_w];
assign c453ibus[temp_w*3 +:temp_w] = v1005obus[temp_w*0 +:temp_w];
assign v1005ibus[data_w*0 +:data_w] = c453obus[data_w*3 +:data_w];
assign c453ibus[temp_w*4 +:temp_w] = v1605obus[temp_w*1 +:temp_w];
assign v1605ibus[data_w*1 +:data_w] = c453obus[data_w*4 +:data_w];
assign c453ibus[temp_w*5 +:temp_w] = v1701obus[temp_w*0 +:temp_w];
assign v1701ibus[data_w*0 +:data_w] = c453obus[data_w*5 +:data_w];
assign c454ibus[temp_w*0 +:temp_w] = v205obus[temp_w*2 +:temp_w];
assign v205ibus[data_w*2 +:data_w] = c454obus[data_w*0 +:data_w];
assign c454ibus[temp_w*1 +:temp_w] = v634obus[temp_w*1 +:temp_w];
assign v634ibus[data_w*1 +:data_w] = c454obus[data_w*1 +:data_w];
assign c454ibus[temp_w*2 +:temp_w] = v879obus[temp_w*2 +:temp_w];
assign v879ibus[data_w*2 +:data_w] = c454obus[data_w*2 +:data_w];
assign c454ibus[temp_w*3 +:temp_w] = v1006obus[temp_w*0 +:temp_w];
assign v1006ibus[data_w*0 +:data_w] = c454obus[data_w*3 +:data_w];
assign c454ibus[temp_w*4 +:temp_w] = v1606obus[temp_w*1 +:temp_w];
assign v1606ibus[data_w*1 +:data_w] = c454obus[data_w*4 +:data_w];
assign c454ibus[temp_w*5 +:temp_w] = v1702obus[temp_w*0 +:temp_w];
assign v1702ibus[data_w*0 +:data_w] = c454obus[data_w*5 +:data_w];
assign c455ibus[temp_w*0 +:temp_w] = v206obus[temp_w*2 +:temp_w];
assign v206ibus[data_w*2 +:data_w] = c455obus[data_w*0 +:data_w];
assign c455ibus[temp_w*1 +:temp_w] = v635obus[temp_w*1 +:temp_w];
assign v635ibus[data_w*1 +:data_w] = c455obus[data_w*1 +:data_w];
assign c455ibus[temp_w*2 +:temp_w] = v880obus[temp_w*2 +:temp_w];
assign v880ibus[data_w*2 +:data_w] = c455obus[data_w*2 +:data_w];
assign c455ibus[temp_w*3 +:temp_w] = v1007obus[temp_w*0 +:temp_w];
assign v1007ibus[data_w*0 +:data_w] = c455obus[data_w*3 +:data_w];
assign c455ibus[temp_w*4 +:temp_w] = v1607obus[temp_w*1 +:temp_w];
assign v1607ibus[data_w*1 +:data_w] = c455obus[data_w*4 +:data_w];
assign c455ibus[temp_w*5 +:temp_w] = v1703obus[temp_w*0 +:temp_w];
assign v1703ibus[data_w*0 +:data_w] = c455obus[data_w*5 +:data_w];
assign c456ibus[temp_w*0 +:temp_w] = v207obus[temp_w*2 +:temp_w];
assign v207ibus[data_w*2 +:data_w] = c456obus[data_w*0 +:data_w];
assign c456ibus[temp_w*1 +:temp_w] = v636obus[temp_w*1 +:temp_w];
assign v636ibus[data_w*1 +:data_w] = c456obus[data_w*1 +:data_w];
assign c456ibus[temp_w*2 +:temp_w] = v881obus[temp_w*2 +:temp_w];
assign v881ibus[data_w*2 +:data_w] = c456obus[data_w*2 +:data_w];
assign c456ibus[temp_w*3 +:temp_w] = v1008obus[temp_w*0 +:temp_w];
assign v1008ibus[data_w*0 +:data_w] = c456obus[data_w*3 +:data_w];
assign c456ibus[temp_w*4 +:temp_w] = v1608obus[temp_w*1 +:temp_w];
assign v1608ibus[data_w*1 +:data_w] = c456obus[data_w*4 +:data_w];
assign c456ibus[temp_w*5 +:temp_w] = v1704obus[temp_w*0 +:temp_w];
assign v1704ibus[data_w*0 +:data_w] = c456obus[data_w*5 +:data_w];
assign c457ibus[temp_w*0 +:temp_w] = v208obus[temp_w*2 +:temp_w];
assign v208ibus[data_w*2 +:data_w] = c457obus[data_w*0 +:data_w];
assign c457ibus[temp_w*1 +:temp_w] = v637obus[temp_w*1 +:temp_w];
assign v637ibus[data_w*1 +:data_w] = c457obus[data_w*1 +:data_w];
assign c457ibus[temp_w*2 +:temp_w] = v882obus[temp_w*2 +:temp_w];
assign v882ibus[data_w*2 +:data_w] = c457obus[data_w*2 +:data_w];
assign c457ibus[temp_w*3 +:temp_w] = v1009obus[temp_w*0 +:temp_w];
assign v1009ibus[data_w*0 +:data_w] = c457obus[data_w*3 +:data_w];
assign c457ibus[temp_w*4 +:temp_w] = v1609obus[temp_w*1 +:temp_w];
assign v1609ibus[data_w*1 +:data_w] = c457obus[data_w*4 +:data_w];
assign c457ibus[temp_w*5 +:temp_w] = v1705obus[temp_w*0 +:temp_w];
assign v1705ibus[data_w*0 +:data_w] = c457obus[data_w*5 +:data_w];
assign c458ibus[temp_w*0 +:temp_w] = v209obus[temp_w*2 +:temp_w];
assign v209ibus[data_w*2 +:data_w] = c458obus[data_w*0 +:data_w];
assign c458ibus[temp_w*1 +:temp_w] = v638obus[temp_w*1 +:temp_w];
assign v638ibus[data_w*1 +:data_w] = c458obus[data_w*1 +:data_w];
assign c458ibus[temp_w*2 +:temp_w] = v883obus[temp_w*2 +:temp_w];
assign v883ibus[data_w*2 +:data_w] = c458obus[data_w*2 +:data_w];
assign c458ibus[temp_w*3 +:temp_w] = v1010obus[temp_w*0 +:temp_w];
assign v1010ibus[data_w*0 +:data_w] = c458obus[data_w*3 +:data_w];
assign c458ibus[temp_w*4 +:temp_w] = v1610obus[temp_w*1 +:temp_w];
assign v1610ibus[data_w*1 +:data_w] = c458obus[data_w*4 +:data_w];
assign c458ibus[temp_w*5 +:temp_w] = v1706obus[temp_w*0 +:temp_w];
assign v1706ibus[data_w*0 +:data_w] = c458obus[data_w*5 +:data_w];
assign c459ibus[temp_w*0 +:temp_w] = v210obus[temp_w*2 +:temp_w];
assign v210ibus[data_w*2 +:data_w] = c459obus[data_w*0 +:data_w];
assign c459ibus[temp_w*1 +:temp_w] = v639obus[temp_w*1 +:temp_w];
assign v639ibus[data_w*1 +:data_w] = c459obus[data_w*1 +:data_w];
assign c459ibus[temp_w*2 +:temp_w] = v884obus[temp_w*2 +:temp_w];
assign v884ibus[data_w*2 +:data_w] = c459obus[data_w*2 +:data_w];
assign c459ibus[temp_w*3 +:temp_w] = v1011obus[temp_w*0 +:temp_w];
assign v1011ibus[data_w*0 +:data_w] = c459obus[data_w*3 +:data_w];
assign c459ibus[temp_w*4 +:temp_w] = v1611obus[temp_w*1 +:temp_w];
assign v1611ibus[data_w*1 +:data_w] = c459obus[data_w*4 +:data_w];
assign c459ibus[temp_w*5 +:temp_w] = v1707obus[temp_w*0 +:temp_w];
assign v1707ibus[data_w*0 +:data_w] = c459obus[data_w*5 +:data_w];
assign c460ibus[temp_w*0 +:temp_w] = v211obus[temp_w*2 +:temp_w];
assign v211ibus[data_w*2 +:data_w] = c460obus[data_w*0 +:data_w];
assign c460ibus[temp_w*1 +:temp_w] = v640obus[temp_w*1 +:temp_w];
assign v640ibus[data_w*1 +:data_w] = c460obus[data_w*1 +:data_w];
assign c460ibus[temp_w*2 +:temp_w] = v885obus[temp_w*2 +:temp_w];
assign v885ibus[data_w*2 +:data_w] = c460obus[data_w*2 +:data_w];
assign c460ibus[temp_w*3 +:temp_w] = v1012obus[temp_w*0 +:temp_w];
assign v1012ibus[data_w*0 +:data_w] = c460obus[data_w*3 +:data_w];
assign c460ibus[temp_w*4 +:temp_w] = v1612obus[temp_w*1 +:temp_w];
assign v1612ibus[data_w*1 +:data_w] = c460obus[data_w*4 +:data_w];
assign c460ibus[temp_w*5 +:temp_w] = v1708obus[temp_w*0 +:temp_w];
assign v1708ibus[data_w*0 +:data_w] = c460obus[data_w*5 +:data_w];
assign c461ibus[temp_w*0 +:temp_w] = v212obus[temp_w*2 +:temp_w];
assign v212ibus[data_w*2 +:data_w] = c461obus[data_w*0 +:data_w];
assign c461ibus[temp_w*1 +:temp_w] = v641obus[temp_w*1 +:temp_w];
assign v641ibus[data_w*1 +:data_w] = c461obus[data_w*1 +:data_w];
assign c461ibus[temp_w*2 +:temp_w] = v886obus[temp_w*2 +:temp_w];
assign v886ibus[data_w*2 +:data_w] = c461obus[data_w*2 +:data_w];
assign c461ibus[temp_w*3 +:temp_w] = v1013obus[temp_w*0 +:temp_w];
assign v1013ibus[data_w*0 +:data_w] = c461obus[data_w*3 +:data_w];
assign c461ibus[temp_w*4 +:temp_w] = v1613obus[temp_w*1 +:temp_w];
assign v1613ibus[data_w*1 +:data_w] = c461obus[data_w*4 +:data_w];
assign c461ibus[temp_w*5 +:temp_w] = v1709obus[temp_w*0 +:temp_w];
assign v1709ibus[data_w*0 +:data_w] = c461obus[data_w*5 +:data_w];
assign c462ibus[temp_w*0 +:temp_w] = v213obus[temp_w*2 +:temp_w];
assign v213ibus[data_w*2 +:data_w] = c462obus[data_w*0 +:data_w];
assign c462ibus[temp_w*1 +:temp_w] = v642obus[temp_w*1 +:temp_w];
assign v642ibus[data_w*1 +:data_w] = c462obus[data_w*1 +:data_w];
assign c462ibus[temp_w*2 +:temp_w] = v887obus[temp_w*2 +:temp_w];
assign v887ibus[data_w*2 +:data_w] = c462obus[data_w*2 +:data_w];
assign c462ibus[temp_w*3 +:temp_w] = v1014obus[temp_w*0 +:temp_w];
assign v1014ibus[data_w*0 +:data_w] = c462obus[data_w*3 +:data_w];
assign c462ibus[temp_w*4 +:temp_w] = v1614obus[temp_w*1 +:temp_w];
assign v1614ibus[data_w*1 +:data_w] = c462obus[data_w*4 +:data_w];
assign c462ibus[temp_w*5 +:temp_w] = v1710obus[temp_w*0 +:temp_w];
assign v1710ibus[data_w*0 +:data_w] = c462obus[data_w*5 +:data_w];
assign c463ibus[temp_w*0 +:temp_w] = v214obus[temp_w*2 +:temp_w];
assign v214ibus[data_w*2 +:data_w] = c463obus[data_w*0 +:data_w];
assign c463ibus[temp_w*1 +:temp_w] = v643obus[temp_w*1 +:temp_w];
assign v643ibus[data_w*1 +:data_w] = c463obus[data_w*1 +:data_w];
assign c463ibus[temp_w*2 +:temp_w] = v888obus[temp_w*2 +:temp_w];
assign v888ibus[data_w*2 +:data_w] = c463obus[data_w*2 +:data_w];
assign c463ibus[temp_w*3 +:temp_w] = v1015obus[temp_w*0 +:temp_w];
assign v1015ibus[data_w*0 +:data_w] = c463obus[data_w*3 +:data_w];
assign c463ibus[temp_w*4 +:temp_w] = v1615obus[temp_w*1 +:temp_w];
assign v1615ibus[data_w*1 +:data_w] = c463obus[data_w*4 +:data_w];
assign c463ibus[temp_w*5 +:temp_w] = v1711obus[temp_w*0 +:temp_w];
assign v1711ibus[data_w*0 +:data_w] = c463obus[data_w*5 +:data_w];
assign c464ibus[temp_w*0 +:temp_w] = v215obus[temp_w*2 +:temp_w];
assign v215ibus[data_w*2 +:data_w] = c464obus[data_w*0 +:data_w];
assign c464ibus[temp_w*1 +:temp_w] = v644obus[temp_w*1 +:temp_w];
assign v644ibus[data_w*1 +:data_w] = c464obus[data_w*1 +:data_w];
assign c464ibus[temp_w*2 +:temp_w] = v889obus[temp_w*2 +:temp_w];
assign v889ibus[data_w*2 +:data_w] = c464obus[data_w*2 +:data_w];
assign c464ibus[temp_w*3 +:temp_w] = v1016obus[temp_w*0 +:temp_w];
assign v1016ibus[data_w*0 +:data_w] = c464obus[data_w*3 +:data_w];
assign c464ibus[temp_w*4 +:temp_w] = v1616obus[temp_w*1 +:temp_w];
assign v1616ibus[data_w*1 +:data_w] = c464obus[data_w*4 +:data_w];
assign c464ibus[temp_w*5 +:temp_w] = v1712obus[temp_w*0 +:temp_w];
assign v1712ibus[data_w*0 +:data_w] = c464obus[data_w*5 +:data_w];
assign c465ibus[temp_w*0 +:temp_w] = v216obus[temp_w*2 +:temp_w];
assign v216ibus[data_w*2 +:data_w] = c465obus[data_w*0 +:data_w];
assign c465ibus[temp_w*1 +:temp_w] = v645obus[temp_w*1 +:temp_w];
assign v645ibus[data_w*1 +:data_w] = c465obus[data_w*1 +:data_w];
assign c465ibus[temp_w*2 +:temp_w] = v890obus[temp_w*2 +:temp_w];
assign v890ibus[data_w*2 +:data_w] = c465obus[data_w*2 +:data_w];
assign c465ibus[temp_w*3 +:temp_w] = v1017obus[temp_w*0 +:temp_w];
assign v1017ibus[data_w*0 +:data_w] = c465obus[data_w*3 +:data_w];
assign c465ibus[temp_w*4 +:temp_w] = v1617obus[temp_w*1 +:temp_w];
assign v1617ibus[data_w*1 +:data_w] = c465obus[data_w*4 +:data_w];
assign c465ibus[temp_w*5 +:temp_w] = v1713obus[temp_w*0 +:temp_w];
assign v1713ibus[data_w*0 +:data_w] = c465obus[data_w*5 +:data_w];
assign c466ibus[temp_w*0 +:temp_w] = v217obus[temp_w*2 +:temp_w];
assign v217ibus[data_w*2 +:data_w] = c466obus[data_w*0 +:data_w];
assign c466ibus[temp_w*1 +:temp_w] = v646obus[temp_w*1 +:temp_w];
assign v646ibus[data_w*1 +:data_w] = c466obus[data_w*1 +:data_w];
assign c466ibus[temp_w*2 +:temp_w] = v891obus[temp_w*2 +:temp_w];
assign v891ibus[data_w*2 +:data_w] = c466obus[data_w*2 +:data_w];
assign c466ibus[temp_w*3 +:temp_w] = v1018obus[temp_w*0 +:temp_w];
assign v1018ibus[data_w*0 +:data_w] = c466obus[data_w*3 +:data_w];
assign c466ibus[temp_w*4 +:temp_w] = v1618obus[temp_w*1 +:temp_w];
assign v1618ibus[data_w*1 +:data_w] = c466obus[data_w*4 +:data_w];
assign c466ibus[temp_w*5 +:temp_w] = v1714obus[temp_w*0 +:temp_w];
assign v1714ibus[data_w*0 +:data_w] = c466obus[data_w*5 +:data_w];
assign c467ibus[temp_w*0 +:temp_w] = v218obus[temp_w*2 +:temp_w];
assign v218ibus[data_w*2 +:data_w] = c467obus[data_w*0 +:data_w];
assign c467ibus[temp_w*1 +:temp_w] = v647obus[temp_w*1 +:temp_w];
assign v647ibus[data_w*1 +:data_w] = c467obus[data_w*1 +:data_w];
assign c467ibus[temp_w*2 +:temp_w] = v892obus[temp_w*2 +:temp_w];
assign v892ibus[data_w*2 +:data_w] = c467obus[data_w*2 +:data_w];
assign c467ibus[temp_w*3 +:temp_w] = v1019obus[temp_w*0 +:temp_w];
assign v1019ibus[data_w*0 +:data_w] = c467obus[data_w*3 +:data_w];
assign c467ibus[temp_w*4 +:temp_w] = v1619obus[temp_w*1 +:temp_w];
assign v1619ibus[data_w*1 +:data_w] = c467obus[data_w*4 +:data_w];
assign c467ibus[temp_w*5 +:temp_w] = v1715obus[temp_w*0 +:temp_w];
assign v1715ibus[data_w*0 +:data_w] = c467obus[data_w*5 +:data_w];
assign c468ibus[temp_w*0 +:temp_w] = v219obus[temp_w*2 +:temp_w];
assign v219ibus[data_w*2 +:data_w] = c468obus[data_w*0 +:data_w];
assign c468ibus[temp_w*1 +:temp_w] = v648obus[temp_w*1 +:temp_w];
assign v648ibus[data_w*1 +:data_w] = c468obus[data_w*1 +:data_w];
assign c468ibus[temp_w*2 +:temp_w] = v893obus[temp_w*2 +:temp_w];
assign v893ibus[data_w*2 +:data_w] = c468obus[data_w*2 +:data_w];
assign c468ibus[temp_w*3 +:temp_w] = v1020obus[temp_w*0 +:temp_w];
assign v1020ibus[data_w*0 +:data_w] = c468obus[data_w*3 +:data_w];
assign c468ibus[temp_w*4 +:temp_w] = v1620obus[temp_w*1 +:temp_w];
assign v1620ibus[data_w*1 +:data_w] = c468obus[data_w*4 +:data_w];
assign c468ibus[temp_w*5 +:temp_w] = v1716obus[temp_w*0 +:temp_w];
assign v1716ibus[data_w*0 +:data_w] = c468obus[data_w*5 +:data_w];
assign c469ibus[temp_w*0 +:temp_w] = v220obus[temp_w*2 +:temp_w];
assign v220ibus[data_w*2 +:data_w] = c469obus[data_w*0 +:data_w];
assign c469ibus[temp_w*1 +:temp_w] = v649obus[temp_w*1 +:temp_w];
assign v649ibus[data_w*1 +:data_w] = c469obus[data_w*1 +:data_w];
assign c469ibus[temp_w*2 +:temp_w] = v894obus[temp_w*2 +:temp_w];
assign v894ibus[data_w*2 +:data_w] = c469obus[data_w*2 +:data_w];
assign c469ibus[temp_w*3 +:temp_w] = v1021obus[temp_w*0 +:temp_w];
assign v1021ibus[data_w*0 +:data_w] = c469obus[data_w*3 +:data_w];
assign c469ibus[temp_w*4 +:temp_w] = v1621obus[temp_w*1 +:temp_w];
assign v1621ibus[data_w*1 +:data_w] = c469obus[data_w*4 +:data_w];
assign c469ibus[temp_w*5 +:temp_w] = v1717obus[temp_w*0 +:temp_w];
assign v1717ibus[data_w*0 +:data_w] = c469obus[data_w*5 +:data_w];
assign c470ibus[temp_w*0 +:temp_w] = v221obus[temp_w*2 +:temp_w];
assign v221ibus[data_w*2 +:data_w] = c470obus[data_w*0 +:data_w];
assign c470ibus[temp_w*1 +:temp_w] = v650obus[temp_w*1 +:temp_w];
assign v650ibus[data_w*1 +:data_w] = c470obus[data_w*1 +:data_w];
assign c470ibus[temp_w*2 +:temp_w] = v895obus[temp_w*2 +:temp_w];
assign v895ibus[data_w*2 +:data_w] = c470obus[data_w*2 +:data_w];
assign c470ibus[temp_w*3 +:temp_w] = v1022obus[temp_w*0 +:temp_w];
assign v1022ibus[data_w*0 +:data_w] = c470obus[data_w*3 +:data_w];
assign c470ibus[temp_w*4 +:temp_w] = v1622obus[temp_w*1 +:temp_w];
assign v1622ibus[data_w*1 +:data_w] = c470obus[data_w*4 +:data_w];
assign c470ibus[temp_w*5 +:temp_w] = v1718obus[temp_w*0 +:temp_w];
assign v1718ibus[data_w*0 +:data_w] = c470obus[data_w*5 +:data_w];
assign c471ibus[temp_w*0 +:temp_w] = v222obus[temp_w*2 +:temp_w];
assign v222ibus[data_w*2 +:data_w] = c471obus[data_w*0 +:data_w];
assign c471ibus[temp_w*1 +:temp_w] = v651obus[temp_w*1 +:temp_w];
assign v651ibus[data_w*1 +:data_w] = c471obus[data_w*1 +:data_w];
assign c471ibus[temp_w*2 +:temp_w] = v896obus[temp_w*2 +:temp_w];
assign v896ibus[data_w*2 +:data_w] = c471obus[data_w*2 +:data_w];
assign c471ibus[temp_w*3 +:temp_w] = v1023obus[temp_w*0 +:temp_w];
assign v1023ibus[data_w*0 +:data_w] = c471obus[data_w*3 +:data_w];
assign c471ibus[temp_w*4 +:temp_w] = v1623obus[temp_w*1 +:temp_w];
assign v1623ibus[data_w*1 +:data_w] = c471obus[data_w*4 +:data_w];
assign c471ibus[temp_w*5 +:temp_w] = v1719obus[temp_w*0 +:temp_w];
assign v1719ibus[data_w*0 +:data_w] = c471obus[data_w*5 +:data_w];
assign c472ibus[temp_w*0 +:temp_w] = v223obus[temp_w*2 +:temp_w];
assign v223ibus[data_w*2 +:data_w] = c472obus[data_w*0 +:data_w];
assign c472ibus[temp_w*1 +:temp_w] = v652obus[temp_w*1 +:temp_w];
assign v652ibus[data_w*1 +:data_w] = c472obus[data_w*1 +:data_w];
assign c472ibus[temp_w*2 +:temp_w] = v897obus[temp_w*2 +:temp_w];
assign v897ibus[data_w*2 +:data_w] = c472obus[data_w*2 +:data_w];
assign c472ibus[temp_w*3 +:temp_w] = v1024obus[temp_w*0 +:temp_w];
assign v1024ibus[data_w*0 +:data_w] = c472obus[data_w*3 +:data_w];
assign c472ibus[temp_w*4 +:temp_w] = v1624obus[temp_w*1 +:temp_w];
assign v1624ibus[data_w*1 +:data_w] = c472obus[data_w*4 +:data_w];
assign c472ibus[temp_w*5 +:temp_w] = v1720obus[temp_w*0 +:temp_w];
assign v1720ibus[data_w*0 +:data_w] = c472obus[data_w*5 +:data_w];
assign c473ibus[temp_w*0 +:temp_w] = v224obus[temp_w*2 +:temp_w];
assign v224ibus[data_w*2 +:data_w] = c473obus[data_w*0 +:data_w];
assign c473ibus[temp_w*1 +:temp_w] = v653obus[temp_w*1 +:temp_w];
assign v653ibus[data_w*1 +:data_w] = c473obus[data_w*1 +:data_w];
assign c473ibus[temp_w*2 +:temp_w] = v898obus[temp_w*2 +:temp_w];
assign v898ibus[data_w*2 +:data_w] = c473obus[data_w*2 +:data_w];
assign c473ibus[temp_w*3 +:temp_w] = v1025obus[temp_w*0 +:temp_w];
assign v1025ibus[data_w*0 +:data_w] = c473obus[data_w*3 +:data_w];
assign c473ibus[temp_w*4 +:temp_w] = v1625obus[temp_w*1 +:temp_w];
assign v1625ibus[data_w*1 +:data_w] = c473obus[data_w*4 +:data_w];
assign c473ibus[temp_w*5 +:temp_w] = v1721obus[temp_w*0 +:temp_w];
assign v1721ibus[data_w*0 +:data_w] = c473obus[data_w*5 +:data_w];
assign c474ibus[temp_w*0 +:temp_w] = v225obus[temp_w*2 +:temp_w];
assign v225ibus[data_w*2 +:data_w] = c474obus[data_w*0 +:data_w];
assign c474ibus[temp_w*1 +:temp_w] = v654obus[temp_w*1 +:temp_w];
assign v654ibus[data_w*1 +:data_w] = c474obus[data_w*1 +:data_w];
assign c474ibus[temp_w*2 +:temp_w] = v899obus[temp_w*2 +:temp_w];
assign v899ibus[data_w*2 +:data_w] = c474obus[data_w*2 +:data_w];
assign c474ibus[temp_w*3 +:temp_w] = v1026obus[temp_w*0 +:temp_w];
assign v1026ibus[data_w*0 +:data_w] = c474obus[data_w*3 +:data_w];
assign c474ibus[temp_w*4 +:temp_w] = v1626obus[temp_w*1 +:temp_w];
assign v1626ibus[data_w*1 +:data_w] = c474obus[data_w*4 +:data_w];
assign c474ibus[temp_w*5 +:temp_w] = v1722obus[temp_w*0 +:temp_w];
assign v1722ibus[data_w*0 +:data_w] = c474obus[data_w*5 +:data_w];
assign c475ibus[temp_w*0 +:temp_w] = v226obus[temp_w*2 +:temp_w];
assign v226ibus[data_w*2 +:data_w] = c475obus[data_w*0 +:data_w];
assign c475ibus[temp_w*1 +:temp_w] = v655obus[temp_w*1 +:temp_w];
assign v655ibus[data_w*1 +:data_w] = c475obus[data_w*1 +:data_w];
assign c475ibus[temp_w*2 +:temp_w] = v900obus[temp_w*2 +:temp_w];
assign v900ibus[data_w*2 +:data_w] = c475obus[data_w*2 +:data_w];
assign c475ibus[temp_w*3 +:temp_w] = v1027obus[temp_w*0 +:temp_w];
assign v1027ibus[data_w*0 +:data_w] = c475obus[data_w*3 +:data_w];
assign c475ibus[temp_w*4 +:temp_w] = v1627obus[temp_w*1 +:temp_w];
assign v1627ibus[data_w*1 +:data_w] = c475obus[data_w*4 +:data_w];
assign c475ibus[temp_w*5 +:temp_w] = v1723obus[temp_w*0 +:temp_w];
assign v1723ibus[data_w*0 +:data_w] = c475obus[data_w*5 +:data_w];
assign c476ibus[temp_w*0 +:temp_w] = v227obus[temp_w*2 +:temp_w];
assign v227ibus[data_w*2 +:data_w] = c476obus[data_w*0 +:data_w];
assign c476ibus[temp_w*1 +:temp_w] = v656obus[temp_w*1 +:temp_w];
assign v656ibus[data_w*1 +:data_w] = c476obus[data_w*1 +:data_w];
assign c476ibus[temp_w*2 +:temp_w] = v901obus[temp_w*2 +:temp_w];
assign v901ibus[data_w*2 +:data_w] = c476obus[data_w*2 +:data_w];
assign c476ibus[temp_w*3 +:temp_w] = v1028obus[temp_w*0 +:temp_w];
assign v1028ibus[data_w*0 +:data_w] = c476obus[data_w*3 +:data_w];
assign c476ibus[temp_w*4 +:temp_w] = v1628obus[temp_w*1 +:temp_w];
assign v1628ibus[data_w*1 +:data_w] = c476obus[data_w*4 +:data_w];
assign c476ibus[temp_w*5 +:temp_w] = v1724obus[temp_w*0 +:temp_w];
assign v1724ibus[data_w*0 +:data_w] = c476obus[data_w*5 +:data_w];
assign c477ibus[temp_w*0 +:temp_w] = v228obus[temp_w*2 +:temp_w];
assign v228ibus[data_w*2 +:data_w] = c477obus[data_w*0 +:data_w];
assign c477ibus[temp_w*1 +:temp_w] = v657obus[temp_w*1 +:temp_w];
assign v657ibus[data_w*1 +:data_w] = c477obus[data_w*1 +:data_w];
assign c477ibus[temp_w*2 +:temp_w] = v902obus[temp_w*2 +:temp_w];
assign v902ibus[data_w*2 +:data_w] = c477obus[data_w*2 +:data_w];
assign c477ibus[temp_w*3 +:temp_w] = v1029obus[temp_w*0 +:temp_w];
assign v1029ibus[data_w*0 +:data_w] = c477obus[data_w*3 +:data_w];
assign c477ibus[temp_w*4 +:temp_w] = v1629obus[temp_w*1 +:temp_w];
assign v1629ibus[data_w*1 +:data_w] = c477obus[data_w*4 +:data_w];
assign c477ibus[temp_w*5 +:temp_w] = v1725obus[temp_w*0 +:temp_w];
assign v1725ibus[data_w*0 +:data_w] = c477obus[data_w*5 +:data_w];
assign c478ibus[temp_w*0 +:temp_w] = v229obus[temp_w*2 +:temp_w];
assign v229ibus[data_w*2 +:data_w] = c478obus[data_w*0 +:data_w];
assign c478ibus[temp_w*1 +:temp_w] = v658obus[temp_w*1 +:temp_w];
assign v658ibus[data_w*1 +:data_w] = c478obus[data_w*1 +:data_w];
assign c478ibus[temp_w*2 +:temp_w] = v903obus[temp_w*2 +:temp_w];
assign v903ibus[data_w*2 +:data_w] = c478obus[data_w*2 +:data_w];
assign c478ibus[temp_w*3 +:temp_w] = v1030obus[temp_w*0 +:temp_w];
assign v1030ibus[data_w*0 +:data_w] = c478obus[data_w*3 +:data_w];
assign c478ibus[temp_w*4 +:temp_w] = v1630obus[temp_w*1 +:temp_w];
assign v1630ibus[data_w*1 +:data_w] = c478obus[data_w*4 +:data_w];
assign c478ibus[temp_w*5 +:temp_w] = v1726obus[temp_w*0 +:temp_w];
assign v1726ibus[data_w*0 +:data_w] = c478obus[data_w*5 +:data_w];
assign c479ibus[temp_w*0 +:temp_w] = v230obus[temp_w*2 +:temp_w];
assign v230ibus[data_w*2 +:data_w] = c479obus[data_w*0 +:data_w];
assign c479ibus[temp_w*1 +:temp_w] = v659obus[temp_w*1 +:temp_w];
assign v659ibus[data_w*1 +:data_w] = c479obus[data_w*1 +:data_w];
assign c479ibus[temp_w*2 +:temp_w] = v904obus[temp_w*2 +:temp_w];
assign v904ibus[data_w*2 +:data_w] = c479obus[data_w*2 +:data_w];
assign c479ibus[temp_w*3 +:temp_w] = v1031obus[temp_w*0 +:temp_w];
assign v1031ibus[data_w*0 +:data_w] = c479obus[data_w*3 +:data_w];
assign c479ibus[temp_w*4 +:temp_w] = v1631obus[temp_w*1 +:temp_w];
assign v1631ibus[data_w*1 +:data_w] = c479obus[data_w*4 +:data_w];
assign c479ibus[temp_w*5 +:temp_w] = v1727obus[temp_w*0 +:temp_w];
assign v1727ibus[data_w*0 +:data_w] = c479obus[data_w*5 +:data_w];
assign c480ibus[temp_w*0 +:temp_w] = v430obus[temp_w*1 +:temp_w];
assign v430ibus[data_w*1 +:data_w] = c480obus[data_w*0 +:data_w];
assign c480ibus[temp_w*1 +:temp_w] = v520obus[temp_w*2 +:temp_w];
assign v520ibus[data_w*2 +:data_w] = c480obus[data_w*1 +:data_w];
assign c480ibus[temp_w*2 +:temp_w] = v754obus[temp_w*2 +:temp_w];
assign v754ibus[data_w*2 +:data_w] = c480obus[data_w*2 +:data_w];
assign c480ibus[temp_w*3 +:temp_w] = v1135obus[temp_w*2 +:temp_w];
assign v1135ibus[data_w*2 +:data_w] = c480obus[data_w*3 +:data_w];
assign c480ibus[temp_w*4 +:temp_w] = v1152obus[temp_w*1 +:temp_w];
assign v1152ibus[data_w*1 +:data_w] = c480obus[data_w*4 +:data_w];
assign c480ibus[temp_w*5 +:temp_w] = v1632obus[temp_w*1 +:temp_w];
assign v1632ibus[data_w*1 +:data_w] = c480obus[data_w*5 +:data_w];
assign c480ibus[temp_w*6 +:temp_w] = v1728obus[temp_w*0 +:temp_w];
assign v1728ibus[data_w*0 +:data_w] = c480obus[data_w*6 +:data_w];
assign c481ibus[temp_w*0 +:temp_w] = v431obus[temp_w*1 +:temp_w];
assign v431ibus[data_w*1 +:data_w] = c481obus[data_w*0 +:data_w];
assign c481ibus[temp_w*1 +:temp_w] = v521obus[temp_w*2 +:temp_w];
assign v521ibus[data_w*2 +:data_w] = c481obus[data_w*1 +:data_w];
assign c481ibus[temp_w*2 +:temp_w] = v755obus[temp_w*2 +:temp_w];
assign v755ibus[data_w*2 +:data_w] = c481obus[data_w*2 +:data_w];
assign c481ibus[temp_w*3 +:temp_w] = v1136obus[temp_w*2 +:temp_w];
assign v1136ibus[data_w*2 +:data_w] = c481obus[data_w*3 +:data_w];
assign c481ibus[temp_w*4 +:temp_w] = v1153obus[temp_w*1 +:temp_w];
assign v1153ibus[data_w*1 +:data_w] = c481obus[data_w*4 +:data_w];
assign c481ibus[temp_w*5 +:temp_w] = v1633obus[temp_w*1 +:temp_w];
assign v1633ibus[data_w*1 +:data_w] = c481obus[data_w*5 +:data_w];
assign c481ibus[temp_w*6 +:temp_w] = v1729obus[temp_w*0 +:temp_w];
assign v1729ibus[data_w*0 +:data_w] = c481obus[data_w*6 +:data_w];
assign c482ibus[temp_w*0 +:temp_w] = v432obus[temp_w*1 +:temp_w];
assign v432ibus[data_w*1 +:data_w] = c482obus[data_w*0 +:data_w];
assign c482ibus[temp_w*1 +:temp_w] = v522obus[temp_w*2 +:temp_w];
assign v522ibus[data_w*2 +:data_w] = c482obus[data_w*1 +:data_w];
assign c482ibus[temp_w*2 +:temp_w] = v756obus[temp_w*2 +:temp_w];
assign v756ibus[data_w*2 +:data_w] = c482obus[data_w*2 +:data_w];
assign c482ibus[temp_w*3 +:temp_w] = v1137obus[temp_w*2 +:temp_w];
assign v1137ibus[data_w*2 +:data_w] = c482obus[data_w*3 +:data_w];
assign c482ibus[temp_w*4 +:temp_w] = v1154obus[temp_w*1 +:temp_w];
assign v1154ibus[data_w*1 +:data_w] = c482obus[data_w*4 +:data_w];
assign c482ibus[temp_w*5 +:temp_w] = v1634obus[temp_w*1 +:temp_w];
assign v1634ibus[data_w*1 +:data_w] = c482obus[data_w*5 +:data_w];
assign c482ibus[temp_w*6 +:temp_w] = v1730obus[temp_w*0 +:temp_w];
assign v1730ibus[data_w*0 +:data_w] = c482obus[data_w*6 +:data_w];
assign c483ibus[temp_w*0 +:temp_w] = v433obus[temp_w*1 +:temp_w];
assign v433ibus[data_w*1 +:data_w] = c483obus[data_w*0 +:data_w];
assign c483ibus[temp_w*1 +:temp_w] = v523obus[temp_w*2 +:temp_w];
assign v523ibus[data_w*2 +:data_w] = c483obus[data_w*1 +:data_w];
assign c483ibus[temp_w*2 +:temp_w] = v757obus[temp_w*2 +:temp_w];
assign v757ibus[data_w*2 +:data_w] = c483obus[data_w*2 +:data_w];
assign c483ibus[temp_w*3 +:temp_w] = v1138obus[temp_w*2 +:temp_w];
assign v1138ibus[data_w*2 +:data_w] = c483obus[data_w*3 +:data_w];
assign c483ibus[temp_w*4 +:temp_w] = v1155obus[temp_w*1 +:temp_w];
assign v1155ibus[data_w*1 +:data_w] = c483obus[data_w*4 +:data_w];
assign c483ibus[temp_w*5 +:temp_w] = v1635obus[temp_w*1 +:temp_w];
assign v1635ibus[data_w*1 +:data_w] = c483obus[data_w*5 +:data_w];
assign c483ibus[temp_w*6 +:temp_w] = v1731obus[temp_w*0 +:temp_w];
assign v1731ibus[data_w*0 +:data_w] = c483obus[data_w*6 +:data_w];
assign c484ibus[temp_w*0 +:temp_w] = v434obus[temp_w*1 +:temp_w];
assign v434ibus[data_w*1 +:data_w] = c484obus[data_w*0 +:data_w];
assign c484ibus[temp_w*1 +:temp_w] = v524obus[temp_w*2 +:temp_w];
assign v524ibus[data_w*2 +:data_w] = c484obus[data_w*1 +:data_w];
assign c484ibus[temp_w*2 +:temp_w] = v758obus[temp_w*2 +:temp_w];
assign v758ibus[data_w*2 +:data_w] = c484obus[data_w*2 +:data_w];
assign c484ibus[temp_w*3 +:temp_w] = v1139obus[temp_w*2 +:temp_w];
assign v1139ibus[data_w*2 +:data_w] = c484obus[data_w*3 +:data_w];
assign c484ibus[temp_w*4 +:temp_w] = v1156obus[temp_w*1 +:temp_w];
assign v1156ibus[data_w*1 +:data_w] = c484obus[data_w*4 +:data_w];
assign c484ibus[temp_w*5 +:temp_w] = v1636obus[temp_w*1 +:temp_w];
assign v1636ibus[data_w*1 +:data_w] = c484obus[data_w*5 +:data_w];
assign c484ibus[temp_w*6 +:temp_w] = v1732obus[temp_w*0 +:temp_w];
assign v1732ibus[data_w*0 +:data_w] = c484obus[data_w*6 +:data_w];
assign c485ibus[temp_w*0 +:temp_w] = v435obus[temp_w*1 +:temp_w];
assign v435ibus[data_w*1 +:data_w] = c485obus[data_w*0 +:data_w];
assign c485ibus[temp_w*1 +:temp_w] = v525obus[temp_w*2 +:temp_w];
assign v525ibus[data_w*2 +:data_w] = c485obus[data_w*1 +:data_w];
assign c485ibus[temp_w*2 +:temp_w] = v759obus[temp_w*2 +:temp_w];
assign v759ibus[data_w*2 +:data_w] = c485obus[data_w*2 +:data_w];
assign c485ibus[temp_w*3 +:temp_w] = v1140obus[temp_w*2 +:temp_w];
assign v1140ibus[data_w*2 +:data_w] = c485obus[data_w*3 +:data_w];
assign c485ibus[temp_w*4 +:temp_w] = v1157obus[temp_w*1 +:temp_w];
assign v1157ibus[data_w*1 +:data_w] = c485obus[data_w*4 +:data_w];
assign c485ibus[temp_w*5 +:temp_w] = v1637obus[temp_w*1 +:temp_w];
assign v1637ibus[data_w*1 +:data_w] = c485obus[data_w*5 +:data_w];
assign c485ibus[temp_w*6 +:temp_w] = v1733obus[temp_w*0 +:temp_w];
assign v1733ibus[data_w*0 +:data_w] = c485obus[data_w*6 +:data_w];
assign c486ibus[temp_w*0 +:temp_w] = v436obus[temp_w*1 +:temp_w];
assign v436ibus[data_w*1 +:data_w] = c486obus[data_w*0 +:data_w];
assign c486ibus[temp_w*1 +:temp_w] = v526obus[temp_w*2 +:temp_w];
assign v526ibus[data_w*2 +:data_w] = c486obus[data_w*1 +:data_w];
assign c486ibus[temp_w*2 +:temp_w] = v760obus[temp_w*2 +:temp_w];
assign v760ibus[data_w*2 +:data_w] = c486obus[data_w*2 +:data_w];
assign c486ibus[temp_w*3 +:temp_w] = v1141obus[temp_w*2 +:temp_w];
assign v1141ibus[data_w*2 +:data_w] = c486obus[data_w*3 +:data_w];
assign c486ibus[temp_w*4 +:temp_w] = v1158obus[temp_w*1 +:temp_w];
assign v1158ibus[data_w*1 +:data_w] = c486obus[data_w*4 +:data_w];
assign c486ibus[temp_w*5 +:temp_w] = v1638obus[temp_w*1 +:temp_w];
assign v1638ibus[data_w*1 +:data_w] = c486obus[data_w*5 +:data_w];
assign c486ibus[temp_w*6 +:temp_w] = v1734obus[temp_w*0 +:temp_w];
assign v1734ibus[data_w*0 +:data_w] = c486obus[data_w*6 +:data_w];
assign c487ibus[temp_w*0 +:temp_w] = v437obus[temp_w*1 +:temp_w];
assign v437ibus[data_w*1 +:data_w] = c487obus[data_w*0 +:data_w];
assign c487ibus[temp_w*1 +:temp_w] = v527obus[temp_w*2 +:temp_w];
assign v527ibus[data_w*2 +:data_w] = c487obus[data_w*1 +:data_w];
assign c487ibus[temp_w*2 +:temp_w] = v761obus[temp_w*2 +:temp_w];
assign v761ibus[data_w*2 +:data_w] = c487obus[data_w*2 +:data_w];
assign c487ibus[temp_w*3 +:temp_w] = v1142obus[temp_w*2 +:temp_w];
assign v1142ibus[data_w*2 +:data_w] = c487obus[data_w*3 +:data_w];
assign c487ibus[temp_w*4 +:temp_w] = v1159obus[temp_w*1 +:temp_w];
assign v1159ibus[data_w*1 +:data_w] = c487obus[data_w*4 +:data_w];
assign c487ibus[temp_w*5 +:temp_w] = v1639obus[temp_w*1 +:temp_w];
assign v1639ibus[data_w*1 +:data_w] = c487obus[data_w*5 +:data_w];
assign c487ibus[temp_w*6 +:temp_w] = v1735obus[temp_w*0 +:temp_w];
assign v1735ibus[data_w*0 +:data_w] = c487obus[data_w*6 +:data_w];
assign c488ibus[temp_w*0 +:temp_w] = v438obus[temp_w*1 +:temp_w];
assign v438ibus[data_w*1 +:data_w] = c488obus[data_w*0 +:data_w];
assign c488ibus[temp_w*1 +:temp_w] = v528obus[temp_w*2 +:temp_w];
assign v528ibus[data_w*2 +:data_w] = c488obus[data_w*1 +:data_w];
assign c488ibus[temp_w*2 +:temp_w] = v762obus[temp_w*2 +:temp_w];
assign v762ibus[data_w*2 +:data_w] = c488obus[data_w*2 +:data_w];
assign c488ibus[temp_w*3 +:temp_w] = v1143obus[temp_w*2 +:temp_w];
assign v1143ibus[data_w*2 +:data_w] = c488obus[data_w*3 +:data_w];
assign c488ibus[temp_w*4 +:temp_w] = v1160obus[temp_w*1 +:temp_w];
assign v1160ibus[data_w*1 +:data_w] = c488obus[data_w*4 +:data_w];
assign c488ibus[temp_w*5 +:temp_w] = v1640obus[temp_w*1 +:temp_w];
assign v1640ibus[data_w*1 +:data_w] = c488obus[data_w*5 +:data_w];
assign c488ibus[temp_w*6 +:temp_w] = v1736obus[temp_w*0 +:temp_w];
assign v1736ibus[data_w*0 +:data_w] = c488obus[data_w*6 +:data_w];
assign c489ibus[temp_w*0 +:temp_w] = v439obus[temp_w*1 +:temp_w];
assign v439ibus[data_w*1 +:data_w] = c489obus[data_w*0 +:data_w];
assign c489ibus[temp_w*1 +:temp_w] = v529obus[temp_w*2 +:temp_w];
assign v529ibus[data_w*2 +:data_w] = c489obus[data_w*1 +:data_w];
assign c489ibus[temp_w*2 +:temp_w] = v763obus[temp_w*2 +:temp_w];
assign v763ibus[data_w*2 +:data_w] = c489obus[data_w*2 +:data_w];
assign c489ibus[temp_w*3 +:temp_w] = v1144obus[temp_w*2 +:temp_w];
assign v1144ibus[data_w*2 +:data_w] = c489obus[data_w*3 +:data_w];
assign c489ibus[temp_w*4 +:temp_w] = v1161obus[temp_w*1 +:temp_w];
assign v1161ibus[data_w*1 +:data_w] = c489obus[data_w*4 +:data_w];
assign c489ibus[temp_w*5 +:temp_w] = v1641obus[temp_w*1 +:temp_w];
assign v1641ibus[data_w*1 +:data_w] = c489obus[data_w*5 +:data_w];
assign c489ibus[temp_w*6 +:temp_w] = v1737obus[temp_w*0 +:temp_w];
assign v1737ibus[data_w*0 +:data_w] = c489obus[data_w*6 +:data_w];
assign c490ibus[temp_w*0 +:temp_w] = v440obus[temp_w*1 +:temp_w];
assign v440ibus[data_w*1 +:data_w] = c490obus[data_w*0 +:data_w];
assign c490ibus[temp_w*1 +:temp_w] = v530obus[temp_w*2 +:temp_w];
assign v530ibus[data_w*2 +:data_w] = c490obus[data_w*1 +:data_w];
assign c490ibus[temp_w*2 +:temp_w] = v764obus[temp_w*2 +:temp_w];
assign v764ibus[data_w*2 +:data_w] = c490obus[data_w*2 +:data_w];
assign c490ibus[temp_w*3 +:temp_w] = v1145obus[temp_w*2 +:temp_w];
assign v1145ibus[data_w*2 +:data_w] = c490obus[data_w*3 +:data_w];
assign c490ibus[temp_w*4 +:temp_w] = v1162obus[temp_w*1 +:temp_w];
assign v1162ibus[data_w*1 +:data_w] = c490obus[data_w*4 +:data_w];
assign c490ibus[temp_w*5 +:temp_w] = v1642obus[temp_w*1 +:temp_w];
assign v1642ibus[data_w*1 +:data_w] = c490obus[data_w*5 +:data_w];
assign c490ibus[temp_w*6 +:temp_w] = v1738obus[temp_w*0 +:temp_w];
assign v1738ibus[data_w*0 +:data_w] = c490obus[data_w*6 +:data_w];
assign c491ibus[temp_w*0 +:temp_w] = v441obus[temp_w*1 +:temp_w];
assign v441ibus[data_w*1 +:data_w] = c491obus[data_w*0 +:data_w];
assign c491ibus[temp_w*1 +:temp_w] = v531obus[temp_w*2 +:temp_w];
assign v531ibus[data_w*2 +:data_w] = c491obus[data_w*1 +:data_w];
assign c491ibus[temp_w*2 +:temp_w] = v765obus[temp_w*2 +:temp_w];
assign v765ibus[data_w*2 +:data_w] = c491obus[data_w*2 +:data_w];
assign c491ibus[temp_w*3 +:temp_w] = v1146obus[temp_w*2 +:temp_w];
assign v1146ibus[data_w*2 +:data_w] = c491obus[data_w*3 +:data_w];
assign c491ibus[temp_w*4 +:temp_w] = v1163obus[temp_w*1 +:temp_w];
assign v1163ibus[data_w*1 +:data_w] = c491obus[data_w*4 +:data_w];
assign c491ibus[temp_w*5 +:temp_w] = v1643obus[temp_w*1 +:temp_w];
assign v1643ibus[data_w*1 +:data_w] = c491obus[data_w*5 +:data_w];
assign c491ibus[temp_w*6 +:temp_w] = v1739obus[temp_w*0 +:temp_w];
assign v1739ibus[data_w*0 +:data_w] = c491obus[data_w*6 +:data_w];
assign c492ibus[temp_w*0 +:temp_w] = v442obus[temp_w*1 +:temp_w];
assign v442ibus[data_w*1 +:data_w] = c492obus[data_w*0 +:data_w];
assign c492ibus[temp_w*1 +:temp_w] = v532obus[temp_w*2 +:temp_w];
assign v532ibus[data_w*2 +:data_w] = c492obus[data_w*1 +:data_w];
assign c492ibus[temp_w*2 +:temp_w] = v766obus[temp_w*2 +:temp_w];
assign v766ibus[data_w*2 +:data_w] = c492obus[data_w*2 +:data_w];
assign c492ibus[temp_w*3 +:temp_w] = v1147obus[temp_w*2 +:temp_w];
assign v1147ibus[data_w*2 +:data_w] = c492obus[data_w*3 +:data_w];
assign c492ibus[temp_w*4 +:temp_w] = v1164obus[temp_w*1 +:temp_w];
assign v1164ibus[data_w*1 +:data_w] = c492obus[data_w*4 +:data_w];
assign c492ibus[temp_w*5 +:temp_w] = v1644obus[temp_w*1 +:temp_w];
assign v1644ibus[data_w*1 +:data_w] = c492obus[data_w*5 +:data_w];
assign c492ibus[temp_w*6 +:temp_w] = v1740obus[temp_w*0 +:temp_w];
assign v1740ibus[data_w*0 +:data_w] = c492obus[data_w*6 +:data_w];
assign c493ibus[temp_w*0 +:temp_w] = v443obus[temp_w*1 +:temp_w];
assign v443ibus[data_w*1 +:data_w] = c493obus[data_w*0 +:data_w];
assign c493ibus[temp_w*1 +:temp_w] = v533obus[temp_w*2 +:temp_w];
assign v533ibus[data_w*2 +:data_w] = c493obus[data_w*1 +:data_w];
assign c493ibus[temp_w*2 +:temp_w] = v767obus[temp_w*2 +:temp_w];
assign v767ibus[data_w*2 +:data_w] = c493obus[data_w*2 +:data_w];
assign c493ibus[temp_w*3 +:temp_w] = v1148obus[temp_w*2 +:temp_w];
assign v1148ibus[data_w*2 +:data_w] = c493obus[data_w*3 +:data_w];
assign c493ibus[temp_w*4 +:temp_w] = v1165obus[temp_w*1 +:temp_w];
assign v1165ibus[data_w*1 +:data_w] = c493obus[data_w*4 +:data_w];
assign c493ibus[temp_w*5 +:temp_w] = v1645obus[temp_w*1 +:temp_w];
assign v1645ibus[data_w*1 +:data_w] = c493obus[data_w*5 +:data_w];
assign c493ibus[temp_w*6 +:temp_w] = v1741obus[temp_w*0 +:temp_w];
assign v1741ibus[data_w*0 +:data_w] = c493obus[data_w*6 +:data_w];
assign c494ibus[temp_w*0 +:temp_w] = v444obus[temp_w*1 +:temp_w];
assign v444ibus[data_w*1 +:data_w] = c494obus[data_w*0 +:data_w];
assign c494ibus[temp_w*1 +:temp_w] = v534obus[temp_w*2 +:temp_w];
assign v534ibus[data_w*2 +:data_w] = c494obus[data_w*1 +:data_w];
assign c494ibus[temp_w*2 +:temp_w] = v672obus[temp_w*2 +:temp_w];
assign v672ibus[data_w*2 +:data_w] = c494obus[data_w*2 +:data_w];
assign c494ibus[temp_w*3 +:temp_w] = v1149obus[temp_w*2 +:temp_w];
assign v1149ibus[data_w*2 +:data_w] = c494obus[data_w*3 +:data_w];
assign c494ibus[temp_w*4 +:temp_w] = v1166obus[temp_w*1 +:temp_w];
assign v1166ibus[data_w*1 +:data_w] = c494obus[data_w*4 +:data_w];
assign c494ibus[temp_w*5 +:temp_w] = v1646obus[temp_w*1 +:temp_w];
assign v1646ibus[data_w*1 +:data_w] = c494obus[data_w*5 +:data_w];
assign c494ibus[temp_w*6 +:temp_w] = v1742obus[temp_w*0 +:temp_w];
assign v1742ibus[data_w*0 +:data_w] = c494obus[data_w*6 +:data_w];
assign c495ibus[temp_w*0 +:temp_w] = v445obus[temp_w*1 +:temp_w];
assign v445ibus[data_w*1 +:data_w] = c495obus[data_w*0 +:data_w];
assign c495ibus[temp_w*1 +:temp_w] = v535obus[temp_w*2 +:temp_w];
assign v535ibus[data_w*2 +:data_w] = c495obus[data_w*1 +:data_w];
assign c495ibus[temp_w*2 +:temp_w] = v673obus[temp_w*2 +:temp_w];
assign v673ibus[data_w*2 +:data_w] = c495obus[data_w*2 +:data_w];
assign c495ibus[temp_w*3 +:temp_w] = v1150obus[temp_w*2 +:temp_w];
assign v1150ibus[data_w*2 +:data_w] = c495obus[data_w*3 +:data_w];
assign c495ibus[temp_w*4 +:temp_w] = v1167obus[temp_w*1 +:temp_w];
assign v1167ibus[data_w*1 +:data_w] = c495obus[data_w*4 +:data_w];
assign c495ibus[temp_w*5 +:temp_w] = v1647obus[temp_w*1 +:temp_w];
assign v1647ibus[data_w*1 +:data_w] = c495obus[data_w*5 +:data_w];
assign c495ibus[temp_w*6 +:temp_w] = v1743obus[temp_w*0 +:temp_w];
assign v1743ibus[data_w*0 +:data_w] = c495obus[data_w*6 +:data_w];
assign c496ibus[temp_w*0 +:temp_w] = v446obus[temp_w*1 +:temp_w];
assign v446ibus[data_w*1 +:data_w] = c496obus[data_w*0 +:data_w];
assign c496ibus[temp_w*1 +:temp_w] = v536obus[temp_w*2 +:temp_w];
assign v536ibus[data_w*2 +:data_w] = c496obus[data_w*1 +:data_w];
assign c496ibus[temp_w*2 +:temp_w] = v674obus[temp_w*2 +:temp_w];
assign v674ibus[data_w*2 +:data_w] = c496obus[data_w*2 +:data_w];
assign c496ibus[temp_w*3 +:temp_w] = v1151obus[temp_w*2 +:temp_w];
assign v1151ibus[data_w*2 +:data_w] = c496obus[data_w*3 +:data_w];
assign c496ibus[temp_w*4 +:temp_w] = v1168obus[temp_w*1 +:temp_w];
assign v1168ibus[data_w*1 +:data_w] = c496obus[data_w*4 +:data_w];
assign c496ibus[temp_w*5 +:temp_w] = v1648obus[temp_w*1 +:temp_w];
assign v1648ibus[data_w*1 +:data_w] = c496obus[data_w*5 +:data_w];
assign c496ibus[temp_w*6 +:temp_w] = v1744obus[temp_w*0 +:temp_w];
assign v1744ibus[data_w*0 +:data_w] = c496obus[data_w*6 +:data_w];
assign c497ibus[temp_w*0 +:temp_w] = v447obus[temp_w*1 +:temp_w];
assign v447ibus[data_w*1 +:data_w] = c497obus[data_w*0 +:data_w];
assign c497ibus[temp_w*1 +:temp_w] = v537obus[temp_w*2 +:temp_w];
assign v537ibus[data_w*2 +:data_w] = c497obus[data_w*1 +:data_w];
assign c497ibus[temp_w*2 +:temp_w] = v675obus[temp_w*2 +:temp_w];
assign v675ibus[data_w*2 +:data_w] = c497obus[data_w*2 +:data_w];
assign c497ibus[temp_w*3 +:temp_w] = v1056obus[temp_w*2 +:temp_w];
assign v1056ibus[data_w*2 +:data_w] = c497obus[data_w*3 +:data_w];
assign c497ibus[temp_w*4 +:temp_w] = v1169obus[temp_w*1 +:temp_w];
assign v1169ibus[data_w*1 +:data_w] = c497obus[data_w*4 +:data_w];
assign c497ibus[temp_w*5 +:temp_w] = v1649obus[temp_w*1 +:temp_w];
assign v1649ibus[data_w*1 +:data_w] = c497obus[data_w*5 +:data_w];
assign c497ibus[temp_w*6 +:temp_w] = v1745obus[temp_w*0 +:temp_w];
assign v1745ibus[data_w*0 +:data_w] = c497obus[data_w*6 +:data_w];
assign c498ibus[temp_w*0 +:temp_w] = v448obus[temp_w*1 +:temp_w];
assign v448ibus[data_w*1 +:data_w] = c498obus[data_w*0 +:data_w];
assign c498ibus[temp_w*1 +:temp_w] = v538obus[temp_w*2 +:temp_w];
assign v538ibus[data_w*2 +:data_w] = c498obus[data_w*1 +:data_w];
assign c498ibus[temp_w*2 +:temp_w] = v676obus[temp_w*2 +:temp_w];
assign v676ibus[data_w*2 +:data_w] = c498obus[data_w*2 +:data_w];
assign c498ibus[temp_w*3 +:temp_w] = v1057obus[temp_w*2 +:temp_w];
assign v1057ibus[data_w*2 +:data_w] = c498obus[data_w*3 +:data_w];
assign c498ibus[temp_w*4 +:temp_w] = v1170obus[temp_w*1 +:temp_w];
assign v1170ibus[data_w*1 +:data_w] = c498obus[data_w*4 +:data_w];
assign c498ibus[temp_w*5 +:temp_w] = v1650obus[temp_w*1 +:temp_w];
assign v1650ibus[data_w*1 +:data_w] = c498obus[data_w*5 +:data_w];
assign c498ibus[temp_w*6 +:temp_w] = v1746obus[temp_w*0 +:temp_w];
assign v1746ibus[data_w*0 +:data_w] = c498obus[data_w*6 +:data_w];
assign c499ibus[temp_w*0 +:temp_w] = v449obus[temp_w*1 +:temp_w];
assign v449ibus[data_w*1 +:data_w] = c499obus[data_w*0 +:data_w];
assign c499ibus[temp_w*1 +:temp_w] = v539obus[temp_w*2 +:temp_w];
assign v539ibus[data_w*2 +:data_w] = c499obus[data_w*1 +:data_w];
assign c499ibus[temp_w*2 +:temp_w] = v677obus[temp_w*2 +:temp_w];
assign v677ibus[data_w*2 +:data_w] = c499obus[data_w*2 +:data_w];
assign c499ibus[temp_w*3 +:temp_w] = v1058obus[temp_w*2 +:temp_w];
assign v1058ibus[data_w*2 +:data_w] = c499obus[data_w*3 +:data_w];
assign c499ibus[temp_w*4 +:temp_w] = v1171obus[temp_w*1 +:temp_w];
assign v1171ibus[data_w*1 +:data_w] = c499obus[data_w*4 +:data_w];
assign c499ibus[temp_w*5 +:temp_w] = v1651obus[temp_w*1 +:temp_w];
assign v1651ibus[data_w*1 +:data_w] = c499obus[data_w*5 +:data_w];
assign c499ibus[temp_w*6 +:temp_w] = v1747obus[temp_w*0 +:temp_w];
assign v1747ibus[data_w*0 +:data_w] = c499obus[data_w*6 +:data_w];
assign c500ibus[temp_w*0 +:temp_w] = v450obus[temp_w*1 +:temp_w];
assign v450ibus[data_w*1 +:data_w] = c500obus[data_w*0 +:data_w];
assign c500ibus[temp_w*1 +:temp_w] = v540obus[temp_w*2 +:temp_w];
assign v540ibus[data_w*2 +:data_w] = c500obus[data_w*1 +:data_w];
assign c500ibus[temp_w*2 +:temp_w] = v678obus[temp_w*2 +:temp_w];
assign v678ibus[data_w*2 +:data_w] = c500obus[data_w*2 +:data_w];
assign c500ibus[temp_w*3 +:temp_w] = v1059obus[temp_w*2 +:temp_w];
assign v1059ibus[data_w*2 +:data_w] = c500obus[data_w*3 +:data_w];
assign c500ibus[temp_w*4 +:temp_w] = v1172obus[temp_w*1 +:temp_w];
assign v1172ibus[data_w*1 +:data_w] = c500obus[data_w*4 +:data_w];
assign c500ibus[temp_w*5 +:temp_w] = v1652obus[temp_w*1 +:temp_w];
assign v1652ibus[data_w*1 +:data_w] = c500obus[data_w*5 +:data_w];
assign c500ibus[temp_w*6 +:temp_w] = v1748obus[temp_w*0 +:temp_w];
assign v1748ibus[data_w*0 +:data_w] = c500obus[data_w*6 +:data_w];
assign c501ibus[temp_w*0 +:temp_w] = v451obus[temp_w*1 +:temp_w];
assign v451ibus[data_w*1 +:data_w] = c501obus[data_w*0 +:data_w];
assign c501ibus[temp_w*1 +:temp_w] = v541obus[temp_w*2 +:temp_w];
assign v541ibus[data_w*2 +:data_w] = c501obus[data_w*1 +:data_w];
assign c501ibus[temp_w*2 +:temp_w] = v679obus[temp_w*2 +:temp_w];
assign v679ibus[data_w*2 +:data_w] = c501obus[data_w*2 +:data_w];
assign c501ibus[temp_w*3 +:temp_w] = v1060obus[temp_w*2 +:temp_w];
assign v1060ibus[data_w*2 +:data_w] = c501obus[data_w*3 +:data_w];
assign c501ibus[temp_w*4 +:temp_w] = v1173obus[temp_w*1 +:temp_w];
assign v1173ibus[data_w*1 +:data_w] = c501obus[data_w*4 +:data_w];
assign c501ibus[temp_w*5 +:temp_w] = v1653obus[temp_w*1 +:temp_w];
assign v1653ibus[data_w*1 +:data_w] = c501obus[data_w*5 +:data_w];
assign c501ibus[temp_w*6 +:temp_w] = v1749obus[temp_w*0 +:temp_w];
assign v1749ibus[data_w*0 +:data_w] = c501obus[data_w*6 +:data_w];
assign c502ibus[temp_w*0 +:temp_w] = v452obus[temp_w*1 +:temp_w];
assign v452ibus[data_w*1 +:data_w] = c502obus[data_w*0 +:data_w];
assign c502ibus[temp_w*1 +:temp_w] = v542obus[temp_w*2 +:temp_w];
assign v542ibus[data_w*2 +:data_w] = c502obus[data_w*1 +:data_w];
assign c502ibus[temp_w*2 +:temp_w] = v680obus[temp_w*2 +:temp_w];
assign v680ibus[data_w*2 +:data_w] = c502obus[data_w*2 +:data_w];
assign c502ibus[temp_w*3 +:temp_w] = v1061obus[temp_w*2 +:temp_w];
assign v1061ibus[data_w*2 +:data_w] = c502obus[data_w*3 +:data_w];
assign c502ibus[temp_w*4 +:temp_w] = v1174obus[temp_w*1 +:temp_w];
assign v1174ibus[data_w*1 +:data_w] = c502obus[data_w*4 +:data_w];
assign c502ibus[temp_w*5 +:temp_w] = v1654obus[temp_w*1 +:temp_w];
assign v1654ibus[data_w*1 +:data_w] = c502obus[data_w*5 +:data_w];
assign c502ibus[temp_w*6 +:temp_w] = v1750obus[temp_w*0 +:temp_w];
assign v1750ibus[data_w*0 +:data_w] = c502obus[data_w*6 +:data_w];
assign c503ibus[temp_w*0 +:temp_w] = v453obus[temp_w*1 +:temp_w];
assign v453ibus[data_w*1 +:data_w] = c503obus[data_w*0 +:data_w];
assign c503ibus[temp_w*1 +:temp_w] = v543obus[temp_w*2 +:temp_w];
assign v543ibus[data_w*2 +:data_w] = c503obus[data_w*1 +:data_w];
assign c503ibus[temp_w*2 +:temp_w] = v681obus[temp_w*2 +:temp_w];
assign v681ibus[data_w*2 +:data_w] = c503obus[data_w*2 +:data_w];
assign c503ibus[temp_w*3 +:temp_w] = v1062obus[temp_w*2 +:temp_w];
assign v1062ibus[data_w*2 +:data_w] = c503obus[data_w*3 +:data_w];
assign c503ibus[temp_w*4 +:temp_w] = v1175obus[temp_w*1 +:temp_w];
assign v1175ibus[data_w*1 +:data_w] = c503obus[data_w*4 +:data_w];
assign c503ibus[temp_w*5 +:temp_w] = v1655obus[temp_w*1 +:temp_w];
assign v1655ibus[data_w*1 +:data_w] = c503obus[data_w*5 +:data_w];
assign c503ibus[temp_w*6 +:temp_w] = v1751obus[temp_w*0 +:temp_w];
assign v1751ibus[data_w*0 +:data_w] = c503obus[data_w*6 +:data_w];
assign c504ibus[temp_w*0 +:temp_w] = v454obus[temp_w*1 +:temp_w];
assign v454ibus[data_w*1 +:data_w] = c504obus[data_w*0 +:data_w];
assign c504ibus[temp_w*1 +:temp_w] = v544obus[temp_w*2 +:temp_w];
assign v544ibus[data_w*2 +:data_w] = c504obus[data_w*1 +:data_w];
assign c504ibus[temp_w*2 +:temp_w] = v682obus[temp_w*2 +:temp_w];
assign v682ibus[data_w*2 +:data_w] = c504obus[data_w*2 +:data_w];
assign c504ibus[temp_w*3 +:temp_w] = v1063obus[temp_w*2 +:temp_w];
assign v1063ibus[data_w*2 +:data_w] = c504obus[data_w*3 +:data_w];
assign c504ibus[temp_w*4 +:temp_w] = v1176obus[temp_w*1 +:temp_w];
assign v1176ibus[data_w*1 +:data_w] = c504obus[data_w*4 +:data_w];
assign c504ibus[temp_w*5 +:temp_w] = v1656obus[temp_w*1 +:temp_w];
assign v1656ibus[data_w*1 +:data_w] = c504obus[data_w*5 +:data_w];
assign c504ibus[temp_w*6 +:temp_w] = v1752obus[temp_w*0 +:temp_w];
assign v1752ibus[data_w*0 +:data_w] = c504obus[data_w*6 +:data_w];
assign c505ibus[temp_w*0 +:temp_w] = v455obus[temp_w*1 +:temp_w];
assign v455ibus[data_w*1 +:data_w] = c505obus[data_w*0 +:data_w];
assign c505ibus[temp_w*1 +:temp_w] = v545obus[temp_w*2 +:temp_w];
assign v545ibus[data_w*2 +:data_w] = c505obus[data_w*1 +:data_w];
assign c505ibus[temp_w*2 +:temp_w] = v683obus[temp_w*2 +:temp_w];
assign v683ibus[data_w*2 +:data_w] = c505obus[data_w*2 +:data_w];
assign c505ibus[temp_w*3 +:temp_w] = v1064obus[temp_w*2 +:temp_w];
assign v1064ibus[data_w*2 +:data_w] = c505obus[data_w*3 +:data_w];
assign c505ibus[temp_w*4 +:temp_w] = v1177obus[temp_w*1 +:temp_w];
assign v1177ibus[data_w*1 +:data_w] = c505obus[data_w*4 +:data_w];
assign c505ibus[temp_w*5 +:temp_w] = v1657obus[temp_w*1 +:temp_w];
assign v1657ibus[data_w*1 +:data_w] = c505obus[data_w*5 +:data_w];
assign c505ibus[temp_w*6 +:temp_w] = v1753obus[temp_w*0 +:temp_w];
assign v1753ibus[data_w*0 +:data_w] = c505obus[data_w*6 +:data_w];
assign c506ibus[temp_w*0 +:temp_w] = v456obus[temp_w*1 +:temp_w];
assign v456ibus[data_w*1 +:data_w] = c506obus[data_w*0 +:data_w];
assign c506ibus[temp_w*1 +:temp_w] = v546obus[temp_w*2 +:temp_w];
assign v546ibus[data_w*2 +:data_w] = c506obus[data_w*1 +:data_w];
assign c506ibus[temp_w*2 +:temp_w] = v684obus[temp_w*2 +:temp_w];
assign v684ibus[data_w*2 +:data_w] = c506obus[data_w*2 +:data_w];
assign c506ibus[temp_w*3 +:temp_w] = v1065obus[temp_w*2 +:temp_w];
assign v1065ibus[data_w*2 +:data_w] = c506obus[data_w*3 +:data_w];
assign c506ibus[temp_w*4 +:temp_w] = v1178obus[temp_w*1 +:temp_w];
assign v1178ibus[data_w*1 +:data_w] = c506obus[data_w*4 +:data_w];
assign c506ibus[temp_w*5 +:temp_w] = v1658obus[temp_w*1 +:temp_w];
assign v1658ibus[data_w*1 +:data_w] = c506obus[data_w*5 +:data_w];
assign c506ibus[temp_w*6 +:temp_w] = v1754obus[temp_w*0 +:temp_w];
assign v1754ibus[data_w*0 +:data_w] = c506obus[data_w*6 +:data_w];
assign c507ibus[temp_w*0 +:temp_w] = v457obus[temp_w*1 +:temp_w];
assign v457ibus[data_w*1 +:data_w] = c507obus[data_w*0 +:data_w];
assign c507ibus[temp_w*1 +:temp_w] = v547obus[temp_w*2 +:temp_w];
assign v547ibus[data_w*2 +:data_w] = c507obus[data_w*1 +:data_w];
assign c507ibus[temp_w*2 +:temp_w] = v685obus[temp_w*2 +:temp_w];
assign v685ibus[data_w*2 +:data_w] = c507obus[data_w*2 +:data_w];
assign c507ibus[temp_w*3 +:temp_w] = v1066obus[temp_w*2 +:temp_w];
assign v1066ibus[data_w*2 +:data_w] = c507obus[data_w*3 +:data_w];
assign c507ibus[temp_w*4 +:temp_w] = v1179obus[temp_w*1 +:temp_w];
assign v1179ibus[data_w*1 +:data_w] = c507obus[data_w*4 +:data_w];
assign c507ibus[temp_w*5 +:temp_w] = v1659obus[temp_w*1 +:temp_w];
assign v1659ibus[data_w*1 +:data_w] = c507obus[data_w*5 +:data_w];
assign c507ibus[temp_w*6 +:temp_w] = v1755obus[temp_w*0 +:temp_w];
assign v1755ibus[data_w*0 +:data_w] = c507obus[data_w*6 +:data_w];
assign c508ibus[temp_w*0 +:temp_w] = v458obus[temp_w*1 +:temp_w];
assign v458ibus[data_w*1 +:data_w] = c508obus[data_w*0 +:data_w];
assign c508ibus[temp_w*1 +:temp_w] = v548obus[temp_w*2 +:temp_w];
assign v548ibus[data_w*2 +:data_w] = c508obus[data_w*1 +:data_w];
assign c508ibus[temp_w*2 +:temp_w] = v686obus[temp_w*2 +:temp_w];
assign v686ibus[data_w*2 +:data_w] = c508obus[data_w*2 +:data_w];
assign c508ibus[temp_w*3 +:temp_w] = v1067obus[temp_w*2 +:temp_w];
assign v1067ibus[data_w*2 +:data_w] = c508obus[data_w*3 +:data_w];
assign c508ibus[temp_w*4 +:temp_w] = v1180obus[temp_w*1 +:temp_w];
assign v1180ibus[data_w*1 +:data_w] = c508obus[data_w*4 +:data_w];
assign c508ibus[temp_w*5 +:temp_w] = v1660obus[temp_w*1 +:temp_w];
assign v1660ibus[data_w*1 +:data_w] = c508obus[data_w*5 +:data_w];
assign c508ibus[temp_w*6 +:temp_w] = v1756obus[temp_w*0 +:temp_w];
assign v1756ibus[data_w*0 +:data_w] = c508obus[data_w*6 +:data_w];
assign c509ibus[temp_w*0 +:temp_w] = v459obus[temp_w*1 +:temp_w];
assign v459ibus[data_w*1 +:data_w] = c509obus[data_w*0 +:data_w];
assign c509ibus[temp_w*1 +:temp_w] = v549obus[temp_w*2 +:temp_w];
assign v549ibus[data_w*2 +:data_w] = c509obus[data_w*1 +:data_w];
assign c509ibus[temp_w*2 +:temp_w] = v687obus[temp_w*2 +:temp_w];
assign v687ibus[data_w*2 +:data_w] = c509obus[data_w*2 +:data_w];
assign c509ibus[temp_w*3 +:temp_w] = v1068obus[temp_w*2 +:temp_w];
assign v1068ibus[data_w*2 +:data_w] = c509obus[data_w*3 +:data_w];
assign c509ibus[temp_w*4 +:temp_w] = v1181obus[temp_w*1 +:temp_w];
assign v1181ibus[data_w*1 +:data_w] = c509obus[data_w*4 +:data_w];
assign c509ibus[temp_w*5 +:temp_w] = v1661obus[temp_w*1 +:temp_w];
assign v1661ibus[data_w*1 +:data_w] = c509obus[data_w*5 +:data_w];
assign c509ibus[temp_w*6 +:temp_w] = v1757obus[temp_w*0 +:temp_w];
assign v1757ibus[data_w*0 +:data_w] = c509obus[data_w*6 +:data_w];
assign c510ibus[temp_w*0 +:temp_w] = v460obus[temp_w*1 +:temp_w];
assign v460ibus[data_w*1 +:data_w] = c510obus[data_w*0 +:data_w];
assign c510ibus[temp_w*1 +:temp_w] = v550obus[temp_w*2 +:temp_w];
assign v550ibus[data_w*2 +:data_w] = c510obus[data_w*1 +:data_w];
assign c510ibus[temp_w*2 +:temp_w] = v688obus[temp_w*2 +:temp_w];
assign v688ibus[data_w*2 +:data_w] = c510obus[data_w*2 +:data_w];
assign c510ibus[temp_w*3 +:temp_w] = v1069obus[temp_w*2 +:temp_w];
assign v1069ibus[data_w*2 +:data_w] = c510obus[data_w*3 +:data_w];
assign c510ibus[temp_w*4 +:temp_w] = v1182obus[temp_w*1 +:temp_w];
assign v1182ibus[data_w*1 +:data_w] = c510obus[data_w*4 +:data_w];
assign c510ibus[temp_w*5 +:temp_w] = v1662obus[temp_w*1 +:temp_w];
assign v1662ibus[data_w*1 +:data_w] = c510obus[data_w*5 +:data_w];
assign c510ibus[temp_w*6 +:temp_w] = v1758obus[temp_w*0 +:temp_w];
assign v1758ibus[data_w*0 +:data_w] = c510obus[data_w*6 +:data_w];
assign c511ibus[temp_w*0 +:temp_w] = v461obus[temp_w*1 +:temp_w];
assign v461ibus[data_w*1 +:data_w] = c511obus[data_w*0 +:data_w];
assign c511ibus[temp_w*1 +:temp_w] = v551obus[temp_w*2 +:temp_w];
assign v551ibus[data_w*2 +:data_w] = c511obus[data_w*1 +:data_w];
assign c511ibus[temp_w*2 +:temp_w] = v689obus[temp_w*2 +:temp_w];
assign v689ibus[data_w*2 +:data_w] = c511obus[data_w*2 +:data_w];
assign c511ibus[temp_w*3 +:temp_w] = v1070obus[temp_w*2 +:temp_w];
assign v1070ibus[data_w*2 +:data_w] = c511obus[data_w*3 +:data_w];
assign c511ibus[temp_w*4 +:temp_w] = v1183obus[temp_w*1 +:temp_w];
assign v1183ibus[data_w*1 +:data_w] = c511obus[data_w*4 +:data_w];
assign c511ibus[temp_w*5 +:temp_w] = v1663obus[temp_w*1 +:temp_w];
assign v1663ibus[data_w*1 +:data_w] = c511obus[data_w*5 +:data_w];
assign c511ibus[temp_w*6 +:temp_w] = v1759obus[temp_w*0 +:temp_w];
assign v1759ibus[data_w*0 +:data_w] = c511obus[data_w*6 +:data_w];
assign c512ibus[temp_w*0 +:temp_w] = v462obus[temp_w*1 +:temp_w];
assign v462ibus[data_w*1 +:data_w] = c512obus[data_w*0 +:data_w];
assign c512ibus[temp_w*1 +:temp_w] = v552obus[temp_w*2 +:temp_w];
assign v552ibus[data_w*2 +:data_w] = c512obus[data_w*1 +:data_w];
assign c512ibus[temp_w*2 +:temp_w] = v690obus[temp_w*2 +:temp_w];
assign v690ibus[data_w*2 +:data_w] = c512obus[data_w*2 +:data_w];
assign c512ibus[temp_w*3 +:temp_w] = v1071obus[temp_w*2 +:temp_w];
assign v1071ibus[data_w*2 +:data_w] = c512obus[data_w*3 +:data_w];
assign c512ibus[temp_w*4 +:temp_w] = v1184obus[temp_w*1 +:temp_w];
assign v1184ibus[data_w*1 +:data_w] = c512obus[data_w*4 +:data_w];
assign c512ibus[temp_w*5 +:temp_w] = v1664obus[temp_w*1 +:temp_w];
assign v1664ibus[data_w*1 +:data_w] = c512obus[data_w*5 +:data_w];
assign c512ibus[temp_w*6 +:temp_w] = v1760obus[temp_w*0 +:temp_w];
assign v1760ibus[data_w*0 +:data_w] = c512obus[data_w*6 +:data_w];
assign c513ibus[temp_w*0 +:temp_w] = v463obus[temp_w*1 +:temp_w];
assign v463ibus[data_w*1 +:data_w] = c513obus[data_w*0 +:data_w];
assign c513ibus[temp_w*1 +:temp_w] = v553obus[temp_w*2 +:temp_w];
assign v553ibus[data_w*2 +:data_w] = c513obus[data_w*1 +:data_w];
assign c513ibus[temp_w*2 +:temp_w] = v691obus[temp_w*2 +:temp_w];
assign v691ibus[data_w*2 +:data_w] = c513obus[data_w*2 +:data_w];
assign c513ibus[temp_w*3 +:temp_w] = v1072obus[temp_w*2 +:temp_w];
assign v1072ibus[data_w*2 +:data_w] = c513obus[data_w*3 +:data_w];
assign c513ibus[temp_w*4 +:temp_w] = v1185obus[temp_w*1 +:temp_w];
assign v1185ibus[data_w*1 +:data_w] = c513obus[data_w*4 +:data_w];
assign c513ibus[temp_w*5 +:temp_w] = v1665obus[temp_w*1 +:temp_w];
assign v1665ibus[data_w*1 +:data_w] = c513obus[data_w*5 +:data_w];
assign c513ibus[temp_w*6 +:temp_w] = v1761obus[temp_w*0 +:temp_w];
assign v1761ibus[data_w*0 +:data_w] = c513obus[data_w*6 +:data_w];
assign c514ibus[temp_w*0 +:temp_w] = v464obus[temp_w*1 +:temp_w];
assign v464ibus[data_w*1 +:data_w] = c514obus[data_w*0 +:data_w];
assign c514ibus[temp_w*1 +:temp_w] = v554obus[temp_w*2 +:temp_w];
assign v554ibus[data_w*2 +:data_w] = c514obus[data_w*1 +:data_w];
assign c514ibus[temp_w*2 +:temp_w] = v692obus[temp_w*2 +:temp_w];
assign v692ibus[data_w*2 +:data_w] = c514obus[data_w*2 +:data_w];
assign c514ibus[temp_w*3 +:temp_w] = v1073obus[temp_w*2 +:temp_w];
assign v1073ibus[data_w*2 +:data_w] = c514obus[data_w*3 +:data_w];
assign c514ibus[temp_w*4 +:temp_w] = v1186obus[temp_w*1 +:temp_w];
assign v1186ibus[data_w*1 +:data_w] = c514obus[data_w*4 +:data_w];
assign c514ibus[temp_w*5 +:temp_w] = v1666obus[temp_w*1 +:temp_w];
assign v1666ibus[data_w*1 +:data_w] = c514obus[data_w*5 +:data_w];
assign c514ibus[temp_w*6 +:temp_w] = v1762obus[temp_w*0 +:temp_w];
assign v1762ibus[data_w*0 +:data_w] = c514obus[data_w*6 +:data_w];
assign c515ibus[temp_w*0 +:temp_w] = v465obus[temp_w*1 +:temp_w];
assign v465ibus[data_w*1 +:data_w] = c515obus[data_w*0 +:data_w];
assign c515ibus[temp_w*1 +:temp_w] = v555obus[temp_w*2 +:temp_w];
assign v555ibus[data_w*2 +:data_w] = c515obus[data_w*1 +:data_w];
assign c515ibus[temp_w*2 +:temp_w] = v693obus[temp_w*2 +:temp_w];
assign v693ibus[data_w*2 +:data_w] = c515obus[data_w*2 +:data_w];
assign c515ibus[temp_w*3 +:temp_w] = v1074obus[temp_w*2 +:temp_w];
assign v1074ibus[data_w*2 +:data_w] = c515obus[data_w*3 +:data_w];
assign c515ibus[temp_w*4 +:temp_w] = v1187obus[temp_w*1 +:temp_w];
assign v1187ibus[data_w*1 +:data_w] = c515obus[data_w*4 +:data_w];
assign c515ibus[temp_w*5 +:temp_w] = v1667obus[temp_w*1 +:temp_w];
assign v1667ibus[data_w*1 +:data_w] = c515obus[data_w*5 +:data_w];
assign c515ibus[temp_w*6 +:temp_w] = v1763obus[temp_w*0 +:temp_w];
assign v1763ibus[data_w*0 +:data_w] = c515obus[data_w*6 +:data_w];
assign c516ibus[temp_w*0 +:temp_w] = v466obus[temp_w*1 +:temp_w];
assign v466ibus[data_w*1 +:data_w] = c516obus[data_w*0 +:data_w];
assign c516ibus[temp_w*1 +:temp_w] = v556obus[temp_w*2 +:temp_w];
assign v556ibus[data_w*2 +:data_w] = c516obus[data_w*1 +:data_w];
assign c516ibus[temp_w*2 +:temp_w] = v694obus[temp_w*2 +:temp_w];
assign v694ibus[data_w*2 +:data_w] = c516obus[data_w*2 +:data_w];
assign c516ibus[temp_w*3 +:temp_w] = v1075obus[temp_w*2 +:temp_w];
assign v1075ibus[data_w*2 +:data_w] = c516obus[data_w*3 +:data_w];
assign c516ibus[temp_w*4 +:temp_w] = v1188obus[temp_w*1 +:temp_w];
assign v1188ibus[data_w*1 +:data_w] = c516obus[data_w*4 +:data_w];
assign c516ibus[temp_w*5 +:temp_w] = v1668obus[temp_w*1 +:temp_w];
assign v1668ibus[data_w*1 +:data_w] = c516obus[data_w*5 +:data_w];
assign c516ibus[temp_w*6 +:temp_w] = v1764obus[temp_w*0 +:temp_w];
assign v1764ibus[data_w*0 +:data_w] = c516obus[data_w*6 +:data_w];
assign c517ibus[temp_w*0 +:temp_w] = v467obus[temp_w*1 +:temp_w];
assign v467ibus[data_w*1 +:data_w] = c517obus[data_w*0 +:data_w];
assign c517ibus[temp_w*1 +:temp_w] = v557obus[temp_w*2 +:temp_w];
assign v557ibus[data_w*2 +:data_w] = c517obus[data_w*1 +:data_w];
assign c517ibus[temp_w*2 +:temp_w] = v695obus[temp_w*2 +:temp_w];
assign v695ibus[data_w*2 +:data_w] = c517obus[data_w*2 +:data_w];
assign c517ibus[temp_w*3 +:temp_w] = v1076obus[temp_w*2 +:temp_w];
assign v1076ibus[data_w*2 +:data_w] = c517obus[data_w*3 +:data_w];
assign c517ibus[temp_w*4 +:temp_w] = v1189obus[temp_w*1 +:temp_w];
assign v1189ibus[data_w*1 +:data_w] = c517obus[data_w*4 +:data_w];
assign c517ibus[temp_w*5 +:temp_w] = v1669obus[temp_w*1 +:temp_w];
assign v1669ibus[data_w*1 +:data_w] = c517obus[data_w*5 +:data_w];
assign c517ibus[temp_w*6 +:temp_w] = v1765obus[temp_w*0 +:temp_w];
assign v1765ibus[data_w*0 +:data_w] = c517obus[data_w*6 +:data_w];
assign c518ibus[temp_w*0 +:temp_w] = v468obus[temp_w*1 +:temp_w];
assign v468ibus[data_w*1 +:data_w] = c518obus[data_w*0 +:data_w];
assign c518ibus[temp_w*1 +:temp_w] = v558obus[temp_w*2 +:temp_w];
assign v558ibus[data_w*2 +:data_w] = c518obus[data_w*1 +:data_w];
assign c518ibus[temp_w*2 +:temp_w] = v696obus[temp_w*2 +:temp_w];
assign v696ibus[data_w*2 +:data_w] = c518obus[data_w*2 +:data_w];
assign c518ibus[temp_w*3 +:temp_w] = v1077obus[temp_w*2 +:temp_w];
assign v1077ibus[data_w*2 +:data_w] = c518obus[data_w*3 +:data_w];
assign c518ibus[temp_w*4 +:temp_w] = v1190obus[temp_w*1 +:temp_w];
assign v1190ibus[data_w*1 +:data_w] = c518obus[data_w*4 +:data_w];
assign c518ibus[temp_w*5 +:temp_w] = v1670obus[temp_w*1 +:temp_w];
assign v1670ibus[data_w*1 +:data_w] = c518obus[data_w*5 +:data_w];
assign c518ibus[temp_w*6 +:temp_w] = v1766obus[temp_w*0 +:temp_w];
assign v1766ibus[data_w*0 +:data_w] = c518obus[data_w*6 +:data_w];
assign c519ibus[temp_w*0 +:temp_w] = v469obus[temp_w*1 +:temp_w];
assign v469ibus[data_w*1 +:data_w] = c519obus[data_w*0 +:data_w];
assign c519ibus[temp_w*1 +:temp_w] = v559obus[temp_w*2 +:temp_w];
assign v559ibus[data_w*2 +:data_w] = c519obus[data_w*1 +:data_w];
assign c519ibus[temp_w*2 +:temp_w] = v697obus[temp_w*2 +:temp_w];
assign v697ibus[data_w*2 +:data_w] = c519obus[data_w*2 +:data_w];
assign c519ibus[temp_w*3 +:temp_w] = v1078obus[temp_w*2 +:temp_w];
assign v1078ibus[data_w*2 +:data_w] = c519obus[data_w*3 +:data_w];
assign c519ibus[temp_w*4 +:temp_w] = v1191obus[temp_w*1 +:temp_w];
assign v1191ibus[data_w*1 +:data_w] = c519obus[data_w*4 +:data_w];
assign c519ibus[temp_w*5 +:temp_w] = v1671obus[temp_w*1 +:temp_w];
assign v1671ibus[data_w*1 +:data_w] = c519obus[data_w*5 +:data_w];
assign c519ibus[temp_w*6 +:temp_w] = v1767obus[temp_w*0 +:temp_w];
assign v1767ibus[data_w*0 +:data_w] = c519obus[data_w*6 +:data_w];
assign c520ibus[temp_w*0 +:temp_w] = v470obus[temp_w*1 +:temp_w];
assign v470ibus[data_w*1 +:data_w] = c520obus[data_w*0 +:data_w];
assign c520ibus[temp_w*1 +:temp_w] = v560obus[temp_w*2 +:temp_w];
assign v560ibus[data_w*2 +:data_w] = c520obus[data_w*1 +:data_w];
assign c520ibus[temp_w*2 +:temp_w] = v698obus[temp_w*2 +:temp_w];
assign v698ibus[data_w*2 +:data_w] = c520obus[data_w*2 +:data_w];
assign c520ibus[temp_w*3 +:temp_w] = v1079obus[temp_w*2 +:temp_w];
assign v1079ibus[data_w*2 +:data_w] = c520obus[data_w*3 +:data_w];
assign c520ibus[temp_w*4 +:temp_w] = v1192obus[temp_w*1 +:temp_w];
assign v1192ibus[data_w*1 +:data_w] = c520obus[data_w*4 +:data_w];
assign c520ibus[temp_w*5 +:temp_w] = v1672obus[temp_w*1 +:temp_w];
assign v1672ibus[data_w*1 +:data_w] = c520obus[data_w*5 +:data_w];
assign c520ibus[temp_w*6 +:temp_w] = v1768obus[temp_w*0 +:temp_w];
assign v1768ibus[data_w*0 +:data_w] = c520obus[data_w*6 +:data_w];
assign c521ibus[temp_w*0 +:temp_w] = v471obus[temp_w*1 +:temp_w];
assign v471ibus[data_w*1 +:data_w] = c521obus[data_w*0 +:data_w];
assign c521ibus[temp_w*1 +:temp_w] = v561obus[temp_w*2 +:temp_w];
assign v561ibus[data_w*2 +:data_w] = c521obus[data_w*1 +:data_w];
assign c521ibus[temp_w*2 +:temp_w] = v699obus[temp_w*2 +:temp_w];
assign v699ibus[data_w*2 +:data_w] = c521obus[data_w*2 +:data_w];
assign c521ibus[temp_w*3 +:temp_w] = v1080obus[temp_w*2 +:temp_w];
assign v1080ibus[data_w*2 +:data_w] = c521obus[data_w*3 +:data_w];
assign c521ibus[temp_w*4 +:temp_w] = v1193obus[temp_w*1 +:temp_w];
assign v1193ibus[data_w*1 +:data_w] = c521obus[data_w*4 +:data_w];
assign c521ibus[temp_w*5 +:temp_w] = v1673obus[temp_w*1 +:temp_w];
assign v1673ibus[data_w*1 +:data_w] = c521obus[data_w*5 +:data_w];
assign c521ibus[temp_w*6 +:temp_w] = v1769obus[temp_w*0 +:temp_w];
assign v1769ibus[data_w*0 +:data_w] = c521obus[data_w*6 +:data_w];
assign c522ibus[temp_w*0 +:temp_w] = v472obus[temp_w*1 +:temp_w];
assign v472ibus[data_w*1 +:data_w] = c522obus[data_w*0 +:data_w];
assign c522ibus[temp_w*1 +:temp_w] = v562obus[temp_w*2 +:temp_w];
assign v562ibus[data_w*2 +:data_w] = c522obus[data_w*1 +:data_w];
assign c522ibus[temp_w*2 +:temp_w] = v700obus[temp_w*2 +:temp_w];
assign v700ibus[data_w*2 +:data_w] = c522obus[data_w*2 +:data_w];
assign c522ibus[temp_w*3 +:temp_w] = v1081obus[temp_w*2 +:temp_w];
assign v1081ibus[data_w*2 +:data_w] = c522obus[data_w*3 +:data_w];
assign c522ibus[temp_w*4 +:temp_w] = v1194obus[temp_w*1 +:temp_w];
assign v1194ibus[data_w*1 +:data_w] = c522obus[data_w*4 +:data_w];
assign c522ibus[temp_w*5 +:temp_w] = v1674obus[temp_w*1 +:temp_w];
assign v1674ibus[data_w*1 +:data_w] = c522obus[data_w*5 +:data_w];
assign c522ibus[temp_w*6 +:temp_w] = v1770obus[temp_w*0 +:temp_w];
assign v1770ibus[data_w*0 +:data_w] = c522obus[data_w*6 +:data_w];
assign c523ibus[temp_w*0 +:temp_w] = v473obus[temp_w*1 +:temp_w];
assign v473ibus[data_w*1 +:data_w] = c523obus[data_w*0 +:data_w];
assign c523ibus[temp_w*1 +:temp_w] = v563obus[temp_w*2 +:temp_w];
assign v563ibus[data_w*2 +:data_w] = c523obus[data_w*1 +:data_w];
assign c523ibus[temp_w*2 +:temp_w] = v701obus[temp_w*2 +:temp_w];
assign v701ibus[data_w*2 +:data_w] = c523obus[data_w*2 +:data_w];
assign c523ibus[temp_w*3 +:temp_w] = v1082obus[temp_w*2 +:temp_w];
assign v1082ibus[data_w*2 +:data_w] = c523obus[data_w*3 +:data_w];
assign c523ibus[temp_w*4 +:temp_w] = v1195obus[temp_w*1 +:temp_w];
assign v1195ibus[data_w*1 +:data_w] = c523obus[data_w*4 +:data_w];
assign c523ibus[temp_w*5 +:temp_w] = v1675obus[temp_w*1 +:temp_w];
assign v1675ibus[data_w*1 +:data_w] = c523obus[data_w*5 +:data_w];
assign c523ibus[temp_w*6 +:temp_w] = v1771obus[temp_w*0 +:temp_w];
assign v1771ibus[data_w*0 +:data_w] = c523obus[data_w*6 +:data_w];
assign c524ibus[temp_w*0 +:temp_w] = v474obus[temp_w*1 +:temp_w];
assign v474ibus[data_w*1 +:data_w] = c524obus[data_w*0 +:data_w];
assign c524ibus[temp_w*1 +:temp_w] = v564obus[temp_w*2 +:temp_w];
assign v564ibus[data_w*2 +:data_w] = c524obus[data_w*1 +:data_w];
assign c524ibus[temp_w*2 +:temp_w] = v702obus[temp_w*2 +:temp_w];
assign v702ibus[data_w*2 +:data_w] = c524obus[data_w*2 +:data_w];
assign c524ibus[temp_w*3 +:temp_w] = v1083obus[temp_w*2 +:temp_w];
assign v1083ibus[data_w*2 +:data_w] = c524obus[data_w*3 +:data_w];
assign c524ibus[temp_w*4 +:temp_w] = v1196obus[temp_w*1 +:temp_w];
assign v1196ibus[data_w*1 +:data_w] = c524obus[data_w*4 +:data_w];
assign c524ibus[temp_w*5 +:temp_w] = v1676obus[temp_w*1 +:temp_w];
assign v1676ibus[data_w*1 +:data_w] = c524obus[data_w*5 +:data_w];
assign c524ibus[temp_w*6 +:temp_w] = v1772obus[temp_w*0 +:temp_w];
assign v1772ibus[data_w*0 +:data_w] = c524obus[data_w*6 +:data_w];
assign c525ibus[temp_w*0 +:temp_w] = v475obus[temp_w*1 +:temp_w];
assign v475ibus[data_w*1 +:data_w] = c525obus[data_w*0 +:data_w];
assign c525ibus[temp_w*1 +:temp_w] = v565obus[temp_w*2 +:temp_w];
assign v565ibus[data_w*2 +:data_w] = c525obus[data_w*1 +:data_w];
assign c525ibus[temp_w*2 +:temp_w] = v703obus[temp_w*2 +:temp_w];
assign v703ibus[data_w*2 +:data_w] = c525obus[data_w*2 +:data_w];
assign c525ibus[temp_w*3 +:temp_w] = v1084obus[temp_w*2 +:temp_w];
assign v1084ibus[data_w*2 +:data_w] = c525obus[data_w*3 +:data_w];
assign c525ibus[temp_w*4 +:temp_w] = v1197obus[temp_w*1 +:temp_w];
assign v1197ibus[data_w*1 +:data_w] = c525obus[data_w*4 +:data_w];
assign c525ibus[temp_w*5 +:temp_w] = v1677obus[temp_w*1 +:temp_w];
assign v1677ibus[data_w*1 +:data_w] = c525obus[data_w*5 +:data_w];
assign c525ibus[temp_w*6 +:temp_w] = v1773obus[temp_w*0 +:temp_w];
assign v1773ibus[data_w*0 +:data_w] = c525obus[data_w*6 +:data_w];
assign c526ibus[temp_w*0 +:temp_w] = v476obus[temp_w*1 +:temp_w];
assign v476ibus[data_w*1 +:data_w] = c526obus[data_w*0 +:data_w];
assign c526ibus[temp_w*1 +:temp_w] = v566obus[temp_w*2 +:temp_w];
assign v566ibus[data_w*2 +:data_w] = c526obus[data_w*1 +:data_w];
assign c526ibus[temp_w*2 +:temp_w] = v704obus[temp_w*2 +:temp_w];
assign v704ibus[data_w*2 +:data_w] = c526obus[data_w*2 +:data_w];
assign c526ibus[temp_w*3 +:temp_w] = v1085obus[temp_w*2 +:temp_w];
assign v1085ibus[data_w*2 +:data_w] = c526obus[data_w*3 +:data_w];
assign c526ibus[temp_w*4 +:temp_w] = v1198obus[temp_w*1 +:temp_w];
assign v1198ibus[data_w*1 +:data_w] = c526obus[data_w*4 +:data_w];
assign c526ibus[temp_w*5 +:temp_w] = v1678obus[temp_w*1 +:temp_w];
assign v1678ibus[data_w*1 +:data_w] = c526obus[data_w*5 +:data_w];
assign c526ibus[temp_w*6 +:temp_w] = v1774obus[temp_w*0 +:temp_w];
assign v1774ibus[data_w*0 +:data_w] = c526obus[data_w*6 +:data_w];
assign c527ibus[temp_w*0 +:temp_w] = v477obus[temp_w*1 +:temp_w];
assign v477ibus[data_w*1 +:data_w] = c527obus[data_w*0 +:data_w];
assign c527ibus[temp_w*1 +:temp_w] = v567obus[temp_w*2 +:temp_w];
assign v567ibus[data_w*2 +:data_w] = c527obus[data_w*1 +:data_w];
assign c527ibus[temp_w*2 +:temp_w] = v705obus[temp_w*2 +:temp_w];
assign v705ibus[data_w*2 +:data_w] = c527obus[data_w*2 +:data_w];
assign c527ibus[temp_w*3 +:temp_w] = v1086obus[temp_w*2 +:temp_w];
assign v1086ibus[data_w*2 +:data_w] = c527obus[data_w*3 +:data_w];
assign c527ibus[temp_w*4 +:temp_w] = v1199obus[temp_w*1 +:temp_w];
assign v1199ibus[data_w*1 +:data_w] = c527obus[data_w*4 +:data_w];
assign c527ibus[temp_w*5 +:temp_w] = v1679obus[temp_w*1 +:temp_w];
assign v1679ibus[data_w*1 +:data_w] = c527obus[data_w*5 +:data_w];
assign c527ibus[temp_w*6 +:temp_w] = v1775obus[temp_w*0 +:temp_w];
assign v1775ibus[data_w*0 +:data_w] = c527obus[data_w*6 +:data_w];
assign c528ibus[temp_w*0 +:temp_w] = v478obus[temp_w*1 +:temp_w];
assign v478ibus[data_w*1 +:data_w] = c528obus[data_w*0 +:data_w];
assign c528ibus[temp_w*1 +:temp_w] = v568obus[temp_w*2 +:temp_w];
assign v568ibus[data_w*2 +:data_w] = c528obus[data_w*1 +:data_w];
assign c528ibus[temp_w*2 +:temp_w] = v706obus[temp_w*2 +:temp_w];
assign v706ibus[data_w*2 +:data_w] = c528obus[data_w*2 +:data_w];
assign c528ibus[temp_w*3 +:temp_w] = v1087obus[temp_w*2 +:temp_w];
assign v1087ibus[data_w*2 +:data_w] = c528obus[data_w*3 +:data_w];
assign c528ibus[temp_w*4 +:temp_w] = v1200obus[temp_w*1 +:temp_w];
assign v1200ibus[data_w*1 +:data_w] = c528obus[data_w*4 +:data_w];
assign c528ibus[temp_w*5 +:temp_w] = v1680obus[temp_w*1 +:temp_w];
assign v1680ibus[data_w*1 +:data_w] = c528obus[data_w*5 +:data_w];
assign c528ibus[temp_w*6 +:temp_w] = v1776obus[temp_w*0 +:temp_w];
assign v1776ibus[data_w*0 +:data_w] = c528obus[data_w*6 +:data_w];
assign c529ibus[temp_w*0 +:temp_w] = v479obus[temp_w*1 +:temp_w];
assign v479ibus[data_w*1 +:data_w] = c529obus[data_w*0 +:data_w];
assign c529ibus[temp_w*1 +:temp_w] = v569obus[temp_w*2 +:temp_w];
assign v569ibus[data_w*2 +:data_w] = c529obus[data_w*1 +:data_w];
assign c529ibus[temp_w*2 +:temp_w] = v707obus[temp_w*2 +:temp_w];
assign v707ibus[data_w*2 +:data_w] = c529obus[data_w*2 +:data_w];
assign c529ibus[temp_w*3 +:temp_w] = v1088obus[temp_w*2 +:temp_w];
assign v1088ibus[data_w*2 +:data_w] = c529obus[data_w*3 +:data_w];
assign c529ibus[temp_w*4 +:temp_w] = v1201obus[temp_w*1 +:temp_w];
assign v1201ibus[data_w*1 +:data_w] = c529obus[data_w*4 +:data_w];
assign c529ibus[temp_w*5 +:temp_w] = v1681obus[temp_w*1 +:temp_w];
assign v1681ibus[data_w*1 +:data_w] = c529obus[data_w*5 +:data_w];
assign c529ibus[temp_w*6 +:temp_w] = v1777obus[temp_w*0 +:temp_w];
assign v1777ibus[data_w*0 +:data_w] = c529obus[data_w*6 +:data_w];
assign c530ibus[temp_w*0 +:temp_w] = v384obus[temp_w*1 +:temp_w];
assign v384ibus[data_w*1 +:data_w] = c530obus[data_w*0 +:data_w];
assign c530ibus[temp_w*1 +:temp_w] = v570obus[temp_w*2 +:temp_w];
assign v570ibus[data_w*2 +:data_w] = c530obus[data_w*1 +:data_w];
assign c530ibus[temp_w*2 +:temp_w] = v708obus[temp_w*2 +:temp_w];
assign v708ibus[data_w*2 +:data_w] = c530obus[data_w*2 +:data_w];
assign c530ibus[temp_w*3 +:temp_w] = v1089obus[temp_w*2 +:temp_w];
assign v1089ibus[data_w*2 +:data_w] = c530obus[data_w*3 +:data_w];
assign c530ibus[temp_w*4 +:temp_w] = v1202obus[temp_w*1 +:temp_w];
assign v1202ibus[data_w*1 +:data_w] = c530obus[data_w*4 +:data_w];
assign c530ibus[temp_w*5 +:temp_w] = v1682obus[temp_w*1 +:temp_w];
assign v1682ibus[data_w*1 +:data_w] = c530obus[data_w*5 +:data_w];
assign c530ibus[temp_w*6 +:temp_w] = v1778obus[temp_w*0 +:temp_w];
assign v1778ibus[data_w*0 +:data_w] = c530obus[data_w*6 +:data_w];
assign c531ibus[temp_w*0 +:temp_w] = v385obus[temp_w*1 +:temp_w];
assign v385ibus[data_w*1 +:data_w] = c531obus[data_w*0 +:data_w];
assign c531ibus[temp_w*1 +:temp_w] = v571obus[temp_w*2 +:temp_w];
assign v571ibus[data_w*2 +:data_w] = c531obus[data_w*1 +:data_w];
assign c531ibus[temp_w*2 +:temp_w] = v709obus[temp_w*2 +:temp_w];
assign v709ibus[data_w*2 +:data_w] = c531obus[data_w*2 +:data_w];
assign c531ibus[temp_w*3 +:temp_w] = v1090obus[temp_w*2 +:temp_w];
assign v1090ibus[data_w*2 +:data_w] = c531obus[data_w*3 +:data_w];
assign c531ibus[temp_w*4 +:temp_w] = v1203obus[temp_w*1 +:temp_w];
assign v1203ibus[data_w*1 +:data_w] = c531obus[data_w*4 +:data_w];
assign c531ibus[temp_w*5 +:temp_w] = v1683obus[temp_w*1 +:temp_w];
assign v1683ibus[data_w*1 +:data_w] = c531obus[data_w*5 +:data_w];
assign c531ibus[temp_w*6 +:temp_w] = v1779obus[temp_w*0 +:temp_w];
assign v1779ibus[data_w*0 +:data_w] = c531obus[data_w*6 +:data_w];
assign c532ibus[temp_w*0 +:temp_w] = v386obus[temp_w*1 +:temp_w];
assign v386ibus[data_w*1 +:data_w] = c532obus[data_w*0 +:data_w];
assign c532ibus[temp_w*1 +:temp_w] = v572obus[temp_w*2 +:temp_w];
assign v572ibus[data_w*2 +:data_w] = c532obus[data_w*1 +:data_w];
assign c532ibus[temp_w*2 +:temp_w] = v710obus[temp_w*2 +:temp_w];
assign v710ibus[data_w*2 +:data_w] = c532obus[data_w*2 +:data_w];
assign c532ibus[temp_w*3 +:temp_w] = v1091obus[temp_w*2 +:temp_w];
assign v1091ibus[data_w*2 +:data_w] = c532obus[data_w*3 +:data_w];
assign c532ibus[temp_w*4 +:temp_w] = v1204obus[temp_w*1 +:temp_w];
assign v1204ibus[data_w*1 +:data_w] = c532obus[data_w*4 +:data_w];
assign c532ibus[temp_w*5 +:temp_w] = v1684obus[temp_w*1 +:temp_w];
assign v1684ibus[data_w*1 +:data_w] = c532obus[data_w*5 +:data_w];
assign c532ibus[temp_w*6 +:temp_w] = v1780obus[temp_w*0 +:temp_w];
assign v1780ibus[data_w*0 +:data_w] = c532obus[data_w*6 +:data_w];
assign c533ibus[temp_w*0 +:temp_w] = v387obus[temp_w*1 +:temp_w];
assign v387ibus[data_w*1 +:data_w] = c533obus[data_w*0 +:data_w];
assign c533ibus[temp_w*1 +:temp_w] = v573obus[temp_w*2 +:temp_w];
assign v573ibus[data_w*2 +:data_w] = c533obus[data_w*1 +:data_w];
assign c533ibus[temp_w*2 +:temp_w] = v711obus[temp_w*2 +:temp_w];
assign v711ibus[data_w*2 +:data_w] = c533obus[data_w*2 +:data_w];
assign c533ibus[temp_w*3 +:temp_w] = v1092obus[temp_w*2 +:temp_w];
assign v1092ibus[data_w*2 +:data_w] = c533obus[data_w*3 +:data_w];
assign c533ibus[temp_w*4 +:temp_w] = v1205obus[temp_w*1 +:temp_w];
assign v1205ibus[data_w*1 +:data_w] = c533obus[data_w*4 +:data_w];
assign c533ibus[temp_w*5 +:temp_w] = v1685obus[temp_w*1 +:temp_w];
assign v1685ibus[data_w*1 +:data_w] = c533obus[data_w*5 +:data_w];
assign c533ibus[temp_w*6 +:temp_w] = v1781obus[temp_w*0 +:temp_w];
assign v1781ibus[data_w*0 +:data_w] = c533obus[data_w*6 +:data_w];
assign c534ibus[temp_w*0 +:temp_w] = v388obus[temp_w*1 +:temp_w];
assign v388ibus[data_w*1 +:data_w] = c534obus[data_w*0 +:data_w];
assign c534ibus[temp_w*1 +:temp_w] = v574obus[temp_w*2 +:temp_w];
assign v574ibus[data_w*2 +:data_w] = c534obus[data_w*1 +:data_w];
assign c534ibus[temp_w*2 +:temp_w] = v712obus[temp_w*2 +:temp_w];
assign v712ibus[data_w*2 +:data_w] = c534obus[data_w*2 +:data_w];
assign c534ibus[temp_w*3 +:temp_w] = v1093obus[temp_w*2 +:temp_w];
assign v1093ibus[data_w*2 +:data_w] = c534obus[data_w*3 +:data_w];
assign c534ibus[temp_w*4 +:temp_w] = v1206obus[temp_w*1 +:temp_w];
assign v1206ibus[data_w*1 +:data_w] = c534obus[data_w*4 +:data_w];
assign c534ibus[temp_w*5 +:temp_w] = v1686obus[temp_w*1 +:temp_w];
assign v1686ibus[data_w*1 +:data_w] = c534obus[data_w*5 +:data_w];
assign c534ibus[temp_w*6 +:temp_w] = v1782obus[temp_w*0 +:temp_w];
assign v1782ibus[data_w*0 +:data_w] = c534obus[data_w*6 +:data_w];
assign c535ibus[temp_w*0 +:temp_w] = v389obus[temp_w*1 +:temp_w];
assign v389ibus[data_w*1 +:data_w] = c535obus[data_w*0 +:data_w];
assign c535ibus[temp_w*1 +:temp_w] = v575obus[temp_w*2 +:temp_w];
assign v575ibus[data_w*2 +:data_w] = c535obus[data_w*1 +:data_w];
assign c535ibus[temp_w*2 +:temp_w] = v713obus[temp_w*2 +:temp_w];
assign v713ibus[data_w*2 +:data_w] = c535obus[data_w*2 +:data_w];
assign c535ibus[temp_w*3 +:temp_w] = v1094obus[temp_w*2 +:temp_w];
assign v1094ibus[data_w*2 +:data_w] = c535obus[data_w*3 +:data_w];
assign c535ibus[temp_w*4 +:temp_w] = v1207obus[temp_w*1 +:temp_w];
assign v1207ibus[data_w*1 +:data_w] = c535obus[data_w*4 +:data_w];
assign c535ibus[temp_w*5 +:temp_w] = v1687obus[temp_w*1 +:temp_w];
assign v1687ibus[data_w*1 +:data_w] = c535obus[data_w*5 +:data_w];
assign c535ibus[temp_w*6 +:temp_w] = v1783obus[temp_w*0 +:temp_w];
assign v1783ibus[data_w*0 +:data_w] = c535obus[data_w*6 +:data_w];
assign c536ibus[temp_w*0 +:temp_w] = v390obus[temp_w*1 +:temp_w];
assign v390ibus[data_w*1 +:data_w] = c536obus[data_w*0 +:data_w];
assign c536ibus[temp_w*1 +:temp_w] = v480obus[temp_w*2 +:temp_w];
assign v480ibus[data_w*2 +:data_w] = c536obus[data_w*1 +:data_w];
assign c536ibus[temp_w*2 +:temp_w] = v714obus[temp_w*2 +:temp_w];
assign v714ibus[data_w*2 +:data_w] = c536obus[data_w*2 +:data_w];
assign c536ibus[temp_w*3 +:temp_w] = v1095obus[temp_w*2 +:temp_w];
assign v1095ibus[data_w*2 +:data_w] = c536obus[data_w*3 +:data_w];
assign c536ibus[temp_w*4 +:temp_w] = v1208obus[temp_w*1 +:temp_w];
assign v1208ibus[data_w*1 +:data_w] = c536obus[data_w*4 +:data_w];
assign c536ibus[temp_w*5 +:temp_w] = v1688obus[temp_w*1 +:temp_w];
assign v1688ibus[data_w*1 +:data_w] = c536obus[data_w*5 +:data_w];
assign c536ibus[temp_w*6 +:temp_w] = v1784obus[temp_w*0 +:temp_w];
assign v1784ibus[data_w*0 +:data_w] = c536obus[data_w*6 +:data_w];
assign c537ibus[temp_w*0 +:temp_w] = v391obus[temp_w*1 +:temp_w];
assign v391ibus[data_w*1 +:data_w] = c537obus[data_w*0 +:data_w];
assign c537ibus[temp_w*1 +:temp_w] = v481obus[temp_w*2 +:temp_w];
assign v481ibus[data_w*2 +:data_w] = c537obus[data_w*1 +:data_w];
assign c537ibus[temp_w*2 +:temp_w] = v715obus[temp_w*2 +:temp_w];
assign v715ibus[data_w*2 +:data_w] = c537obus[data_w*2 +:data_w];
assign c537ibus[temp_w*3 +:temp_w] = v1096obus[temp_w*2 +:temp_w];
assign v1096ibus[data_w*2 +:data_w] = c537obus[data_w*3 +:data_w];
assign c537ibus[temp_w*4 +:temp_w] = v1209obus[temp_w*1 +:temp_w];
assign v1209ibus[data_w*1 +:data_w] = c537obus[data_w*4 +:data_w];
assign c537ibus[temp_w*5 +:temp_w] = v1689obus[temp_w*1 +:temp_w];
assign v1689ibus[data_w*1 +:data_w] = c537obus[data_w*5 +:data_w];
assign c537ibus[temp_w*6 +:temp_w] = v1785obus[temp_w*0 +:temp_w];
assign v1785ibus[data_w*0 +:data_w] = c537obus[data_w*6 +:data_w];
assign c538ibus[temp_w*0 +:temp_w] = v392obus[temp_w*1 +:temp_w];
assign v392ibus[data_w*1 +:data_w] = c538obus[data_w*0 +:data_w];
assign c538ibus[temp_w*1 +:temp_w] = v482obus[temp_w*2 +:temp_w];
assign v482ibus[data_w*2 +:data_w] = c538obus[data_w*1 +:data_w];
assign c538ibus[temp_w*2 +:temp_w] = v716obus[temp_w*2 +:temp_w];
assign v716ibus[data_w*2 +:data_w] = c538obus[data_w*2 +:data_w];
assign c538ibus[temp_w*3 +:temp_w] = v1097obus[temp_w*2 +:temp_w];
assign v1097ibus[data_w*2 +:data_w] = c538obus[data_w*3 +:data_w];
assign c538ibus[temp_w*4 +:temp_w] = v1210obus[temp_w*1 +:temp_w];
assign v1210ibus[data_w*1 +:data_w] = c538obus[data_w*4 +:data_w];
assign c538ibus[temp_w*5 +:temp_w] = v1690obus[temp_w*1 +:temp_w];
assign v1690ibus[data_w*1 +:data_w] = c538obus[data_w*5 +:data_w];
assign c538ibus[temp_w*6 +:temp_w] = v1786obus[temp_w*0 +:temp_w];
assign v1786ibus[data_w*0 +:data_w] = c538obus[data_w*6 +:data_w];
assign c539ibus[temp_w*0 +:temp_w] = v393obus[temp_w*1 +:temp_w];
assign v393ibus[data_w*1 +:data_w] = c539obus[data_w*0 +:data_w];
assign c539ibus[temp_w*1 +:temp_w] = v483obus[temp_w*2 +:temp_w];
assign v483ibus[data_w*2 +:data_w] = c539obus[data_w*1 +:data_w];
assign c539ibus[temp_w*2 +:temp_w] = v717obus[temp_w*2 +:temp_w];
assign v717ibus[data_w*2 +:data_w] = c539obus[data_w*2 +:data_w];
assign c539ibus[temp_w*3 +:temp_w] = v1098obus[temp_w*2 +:temp_w];
assign v1098ibus[data_w*2 +:data_w] = c539obus[data_w*3 +:data_w];
assign c539ibus[temp_w*4 +:temp_w] = v1211obus[temp_w*1 +:temp_w];
assign v1211ibus[data_w*1 +:data_w] = c539obus[data_w*4 +:data_w];
assign c539ibus[temp_w*5 +:temp_w] = v1691obus[temp_w*1 +:temp_w];
assign v1691ibus[data_w*1 +:data_w] = c539obus[data_w*5 +:data_w];
assign c539ibus[temp_w*6 +:temp_w] = v1787obus[temp_w*0 +:temp_w];
assign v1787ibus[data_w*0 +:data_w] = c539obus[data_w*6 +:data_w];
assign c540ibus[temp_w*0 +:temp_w] = v394obus[temp_w*1 +:temp_w];
assign v394ibus[data_w*1 +:data_w] = c540obus[data_w*0 +:data_w];
assign c540ibus[temp_w*1 +:temp_w] = v484obus[temp_w*2 +:temp_w];
assign v484ibus[data_w*2 +:data_w] = c540obus[data_w*1 +:data_w];
assign c540ibus[temp_w*2 +:temp_w] = v718obus[temp_w*2 +:temp_w];
assign v718ibus[data_w*2 +:data_w] = c540obus[data_w*2 +:data_w];
assign c540ibus[temp_w*3 +:temp_w] = v1099obus[temp_w*2 +:temp_w];
assign v1099ibus[data_w*2 +:data_w] = c540obus[data_w*3 +:data_w];
assign c540ibus[temp_w*4 +:temp_w] = v1212obus[temp_w*1 +:temp_w];
assign v1212ibus[data_w*1 +:data_w] = c540obus[data_w*4 +:data_w];
assign c540ibus[temp_w*5 +:temp_w] = v1692obus[temp_w*1 +:temp_w];
assign v1692ibus[data_w*1 +:data_w] = c540obus[data_w*5 +:data_w];
assign c540ibus[temp_w*6 +:temp_w] = v1788obus[temp_w*0 +:temp_w];
assign v1788ibus[data_w*0 +:data_w] = c540obus[data_w*6 +:data_w];
assign c541ibus[temp_w*0 +:temp_w] = v395obus[temp_w*1 +:temp_w];
assign v395ibus[data_w*1 +:data_w] = c541obus[data_w*0 +:data_w];
assign c541ibus[temp_w*1 +:temp_w] = v485obus[temp_w*2 +:temp_w];
assign v485ibus[data_w*2 +:data_w] = c541obus[data_w*1 +:data_w];
assign c541ibus[temp_w*2 +:temp_w] = v719obus[temp_w*2 +:temp_w];
assign v719ibus[data_w*2 +:data_w] = c541obus[data_w*2 +:data_w];
assign c541ibus[temp_w*3 +:temp_w] = v1100obus[temp_w*2 +:temp_w];
assign v1100ibus[data_w*2 +:data_w] = c541obus[data_w*3 +:data_w];
assign c541ibus[temp_w*4 +:temp_w] = v1213obus[temp_w*1 +:temp_w];
assign v1213ibus[data_w*1 +:data_w] = c541obus[data_w*4 +:data_w];
assign c541ibus[temp_w*5 +:temp_w] = v1693obus[temp_w*1 +:temp_w];
assign v1693ibus[data_w*1 +:data_w] = c541obus[data_w*5 +:data_w];
assign c541ibus[temp_w*6 +:temp_w] = v1789obus[temp_w*0 +:temp_w];
assign v1789ibus[data_w*0 +:data_w] = c541obus[data_w*6 +:data_w];
assign c542ibus[temp_w*0 +:temp_w] = v396obus[temp_w*1 +:temp_w];
assign v396ibus[data_w*1 +:data_w] = c542obus[data_w*0 +:data_w];
assign c542ibus[temp_w*1 +:temp_w] = v486obus[temp_w*2 +:temp_w];
assign v486ibus[data_w*2 +:data_w] = c542obus[data_w*1 +:data_w];
assign c542ibus[temp_w*2 +:temp_w] = v720obus[temp_w*2 +:temp_w];
assign v720ibus[data_w*2 +:data_w] = c542obus[data_w*2 +:data_w];
assign c542ibus[temp_w*3 +:temp_w] = v1101obus[temp_w*2 +:temp_w];
assign v1101ibus[data_w*2 +:data_w] = c542obus[data_w*3 +:data_w];
assign c542ibus[temp_w*4 +:temp_w] = v1214obus[temp_w*1 +:temp_w];
assign v1214ibus[data_w*1 +:data_w] = c542obus[data_w*4 +:data_w];
assign c542ibus[temp_w*5 +:temp_w] = v1694obus[temp_w*1 +:temp_w];
assign v1694ibus[data_w*1 +:data_w] = c542obus[data_w*5 +:data_w];
assign c542ibus[temp_w*6 +:temp_w] = v1790obus[temp_w*0 +:temp_w];
assign v1790ibus[data_w*0 +:data_w] = c542obus[data_w*6 +:data_w];
assign c543ibus[temp_w*0 +:temp_w] = v397obus[temp_w*1 +:temp_w];
assign v397ibus[data_w*1 +:data_w] = c543obus[data_w*0 +:data_w];
assign c543ibus[temp_w*1 +:temp_w] = v487obus[temp_w*2 +:temp_w];
assign v487ibus[data_w*2 +:data_w] = c543obus[data_w*1 +:data_w];
assign c543ibus[temp_w*2 +:temp_w] = v721obus[temp_w*2 +:temp_w];
assign v721ibus[data_w*2 +:data_w] = c543obus[data_w*2 +:data_w];
assign c543ibus[temp_w*3 +:temp_w] = v1102obus[temp_w*2 +:temp_w];
assign v1102ibus[data_w*2 +:data_w] = c543obus[data_w*3 +:data_w];
assign c543ibus[temp_w*4 +:temp_w] = v1215obus[temp_w*1 +:temp_w];
assign v1215ibus[data_w*1 +:data_w] = c543obus[data_w*4 +:data_w];
assign c543ibus[temp_w*5 +:temp_w] = v1695obus[temp_w*1 +:temp_w];
assign v1695ibus[data_w*1 +:data_w] = c543obus[data_w*5 +:data_w];
assign c543ibus[temp_w*6 +:temp_w] = v1791obus[temp_w*0 +:temp_w];
assign v1791ibus[data_w*0 +:data_w] = c543obus[data_w*6 +:data_w];
assign c544ibus[temp_w*0 +:temp_w] = v398obus[temp_w*1 +:temp_w];
assign v398ibus[data_w*1 +:data_w] = c544obus[data_w*0 +:data_w];
assign c544ibus[temp_w*1 +:temp_w] = v488obus[temp_w*2 +:temp_w];
assign v488ibus[data_w*2 +:data_w] = c544obus[data_w*1 +:data_w];
assign c544ibus[temp_w*2 +:temp_w] = v722obus[temp_w*2 +:temp_w];
assign v722ibus[data_w*2 +:data_w] = c544obus[data_w*2 +:data_w];
assign c544ibus[temp_w*3 +:temp_w] = v1103obus[temp_w*2 +:temp_w];
assign v1103ibus[data_w*2 +:data_w] = c544obus[data_w*3 +:data_w];
assign c544ibus[temp_w*4 +:temp_w] = v1216obus[temp_w*1 +:temp_w];
assign v1216ibus[data_w*1 +:data_w] = c544obus[data_w*4 +:data_w];
assign c544ibus[temp_w*5 +:temp_w] = v1696obus[temp_w*1 +:temp_w];
assign v1696ibus[data_w*1 +:data_w] = c544obus[data_w*5 +:data_w];
assign c544ibus[temp_w*6 +:temp_w] = v1792obus[temp_w*0 +:temp_w];
assign v1792ibus[data_w*0 +:data_w] = c544obus[data_w*6 +:data_w];
assign c545ibus[temp_w*0 +:temp_w] = v399obus[temp_w*1 +:temp_w];
assign v399ibus[data_w*1 +:data_w] = c545obus[data_w*0 +:data_w];
assign c545ibus[temp_w*1 +:temp_w] = v489obus[temp_w*2 +:temp_w];
assign v489ibus[data_w*2 +:data_w] = c545obus[data_w*1 +:data_w];
assign c545ibus[temp_w*2 +:temp_w] = v723obus[temp_w*2 +:temp_w];
assign v723ibus[data_w*2 +:data_w] = c545obus[data_w*2 +:data_w];
assign c545ibus[temp_w*3 +:temp_w] = v1104obus[temp_w*2 +:temp_w];
assign v1104ibus[data_w*2 +:data_w] = c545obus[data_w*3 +:data_w];
assign c545ibus[temp_w*4 +:temp_w] = v1217obus[temp_w*1 +:temp_w];
assign v1217ibus[data_w*1 +:data_w] = c545obus[data_w*4 +:data_w];
assign c545ibus[temp_w*5 +:temp_w] = v1697obus[temp_w*1 +:temp_w];
assign v1697ibus[data_w*1 +:data_w] = c545obus[data_w*5 +:data_w];
assign c545ibus[temp_w*6 +:temp_w] = v1793obus[temp_w*0 +:temp_w];
assign v1793ibus[data_w*0 +:data_w] = c545obus[data_w*6 +:data_w];
assign c546ibus[temp_w*0 +:temp_w] = v400obus[temp_w*1 +:temp_w];
assign v400ibus[data_w*1 +:data_w] = c546obus[data_w*0 +:data_w];
assign c546ibus[temp_w*1 +:temp_w] = v490obus[temp_w*2 +:temp_w];
assign v490ibus[data_w*2 +:data_w] = c546obus[data_w*1 +:data_w];
assign c546ibus[temp_w*2 +:temp_w] = v724obus[temp_w*2 +:temp_w];
assign v724ibus[data_w*2 +:data_w] = c546obus[data_w*2 +:data_w];
assign c546ibus[temp_w*3 +:temp_w] = v1105obus[temp_w*2 +:temp_w];
assign v1105ibus[data_w*2 +:data_w] = c546obus[data_w*3 +:data_w];
assign c546ibus[temp_w*4 +:temp_w] = v1218obus[temp_w*1 +:temp_w];
assign v1218ibus[data_w*1 +:data_w] = c546obus[data_w*4 +:data_w];
assign c546ibus[temp_w*5 +:temp_w] = v1698obus[temp_w*1 +:temp_w];
assign v1698ibus[data_w*1 +:data_w] = c546obus[data_w*5 +:data_w];
assign c546ibus[temp_w*6 +:temp_w] = v1794obus[temp_w*0 +:temp_w];
assign v1794ibus[data_w*0 +:data_w] = c546obus[data_w*6 +:data_w];
assign c547ibus[temp_w*0 +:temp_w] = v401obus[temp_w*1 +:temp_w];
assign v401ibus[data_w*1 +:data_w] = c547obus[data_w*0 +:data_w];
assign c547ibus[temp_w*1 +:temp_w] = v491obus[temp_w*2 +:temp_w];
assign v491ibus[data_w*2 +:data_w] = c547obus[data_w*1 +:data_w];
assign c547ibus[temp_w*2 +:temp_w] = v725obus[temp_w*2 +:temp_w];
assign v725ibus[data_w*2 +:data_w] = c547obus[data_w*2 +:data_w];
assign c547ibus[temp_w*3 +:temp_w] = v1106obus[temp_w*2 +:temp_w];
assign v1106ibus[data_w*2 +:data_w] = c547obus[data_w*3 +:data_w];
assign c547ibus[temp_w*4 +:temp_w] = v1219obus[temp_w*1 +:temp_w];
assign v1219ibus[data_w*1 +:data_w] = c547obus[data_w*4 +:data_w];
assign c547ibus[temp_w*5 +:temp_w] = v1699obus[temp_w*1 +:temp_w];
assign v1699ibus[data_w*1 +:data_w] = c547obus[data_w*5 +:data_w];
assign c547ibus[temp_w*6 +:temp_w] = v1795obus[temp_w*0 +:temp_w];
assign v1795ibus[data_w*0 +:data_w] = c547obus[data_w*6 +:data_w];
assign c548ibus[temp_w*0 +:temp_w] = v402obus[temp_w*1 +:temp_w];
assign v402ibus[data_w*1 +:data_w] = c548obus[data_w*0 +:data_w];
assign c548ibus[temp_w*1 +:temp_w] = v492obus[temp_w*2 +:temp_w];
assign v492ibus[data_w*2 +:data_w] = c548obus[data_w*1 +:data_w];
assign c548ibus[temp_w*2 +:temp_w] = v726obus[temp_w*2 +:temp_w];
assign v726ibus[data_w*2 +:data_w] = c548obus[data_w*2 +:data_w];
assign c548ibus[temp_w*3 +:temp_w] = v1107obus[temp_w*2 +:temp_w];
assign v1107ibus[data_w*2 +:data_w] = c548obus[data_w*3 +:data_w];
assign c548ibus[temp_w*4 +:temp_w] = v1220obus[temp_w*1 +:temp_w];
assign v1220ibus[data_w*1 +:data_w] = c548obus[data_w*4 +:data_w];
assign c548ibus[temp_w*5 +:temp_w] = v1700obus[temp_w*1 +:temp_w];
assign v1700ibus[data_w*1 +:data_w] = c548obus[data_w*5 +:data_w];
assign c548ibus[temp_w*6 +:temp_w] = v1796obus[temp_w*0 +:temp_w];
assign v1796ibus[data_w*0 +:data_w] = c548obus[data_w*6 +:data_w];
assign c549ibus[temp_w*0 +:temp_w] = v403obus[temp_w*1 +:temp_w];
assign v403ibus[data_w*1 +:data_w] = c549obus[data_w*0 +:data_w];
assign c549ibus[temp_w*1 +:temp_w] = v493obus[temp_w*2 +:temp_w];
assign v493ibus[data_w*2 +:data_w] = c549obus[data_w*1 +:data_w];
assign c549ibus[temp_w*2 +:temp_w] = v727obus[temp_w*2 +:temp_w];
assign v727ibus[data_w*2 +:data_w] = c549obus[data_w*2 +:data_w];
assign c549ibus[temp_w*3 +:temp_w] = v1108obus[temp_w*2 +:temp_w];
assign v1108ibus[data_w*2 +:data_w] = c549obus[data_w*3 +:data_w];
assign c549ibus[temp_w*4 +:temp_w] = v1221obus[temp_w*1 +:temp_w];
assign v1221ibus[data_w*1 +:data_w] = c549obus[data_w*4 +:data_w];
assign c549ibus[temp_w*5 +:temp_w] = v1701obus[temp_w*1 +:temp_w];
assign v1701ibus[data_w*1 +:data_w] = c549obus[data_w*5 +:data_w];
assign c549ibus[temp_w*6 +:temp_w] = v1797obus[temp_w*0 +:temp_w];
assign v1797ibus[data_w*0 +:data_w] = c549obus[data_w*6 +:data_w];
assign c550ibus[temp_w*0 +:temp_w] = v404obus[temp_w*1 +:temp_w];
assign v404ibus[data_w*1 +:data_w] = c550obus[data_w*0 +:data_w];
assign c550ibus[temp_w*1 +:temp_w] = v494obus[temp_w*2 +:temp_w];
assign v494ibus[data_w*2 +:data_w] = c550obus[data_w*1 +:data_w];
assign c550ibus[temp_w*2 +:temp_w] = v728obus[temp_w*2 +:temp_w];
assign v728ibus[data_w*2 +:data_w] = c550obus[data_w*2 +:data_w];
assign c550ibus[temp_w*3 +:temp_w] = v1109obus[temp_w*2 +:temp_w];
assign v1109ibus[data_w*2 +:data_w] = c550obus[data_w*3 +:data_w];
assign c550ibus[temp_w*4 +:temp_w] = v1222obus[temp_w*1 +:temp_w];
assign v1222ibus[data_w*1 +:data_w] = c550obus[data_w*4 +:data_w];
assign c550ibus[temp_w*5 +:temp_w] = v1702obus[temp_w*1 +:temp_w];
assign v1702ibus[data_w*1 +:data_w] = c550obus[data_w*5 +:data_w];
assign c550ibus[temp_w*6 +:temp_w] = v1798obus[temp_w*0 +:temp_w];
assign v1798ibus[data_w*0 +:data_w] = c550obus[data_w*6 +:data_w];
assign c551ibus[temp_w*0 +:temp_w] = v405obus[temp_w*1 +:temp_w];
assign v405ibus[data_w*1 +:data_w] = c551obus[data_w*0 +:data_w];
assign c551ibus[temp_w*1 +:temp_w] = v495obus[temp_w*2 +:temp_w];
assign v495ibus[data_w*2 +:data_w] = c551obus[data_w*1 +:data_w];
assign c551ibus[temp_w*2 +:temp_w] = v729obus[temp_w*2 +:temp_w];
assign v729ibus[data_w*2 +:data_w] = c551obus[data_w*2 +:data_w];
assign c551ibus[temp_w*3 +:temp_w] = v1110obus[temp_w*2 +:temp_w];
assign v1110ibus[data_w*2 +:data_w] = c551obus[data_w*3 +:data_w];
assign c551ibus[temp_w*4 +:temp_w] = v1223obus[temp_w*1 +:temp_w];
assign v1223ibus[data_w*1 +:data_w] = c551obus[data_w*4 +:data_w];
assign c551ibus[temp_w*5 +:temp_w] = v1703obus[temp_w*1 +:temp_w];
assign v1703ibus[data_w*1 +:data_w] = c551obus[data_w*5 +:data_w];
assign c551ibus[temp_w*6 +:temp_w] = v1799obus[temp_w*0 +:temp_w];
assign v1799ibus[data_w*0 +:data_w] = c551obus[data_w*6 +:data_w];
assign c552ibus[temp_w*0 +:temp_w] = v406obus[temp_w*1 +:temp_w];
assign v406ibus[data_w*1 +:data_w] = c552obus[data_w*0 +:data_w];
assign c552ibus[temp_w*1 +:temp_w] = v496obus[temp_w*2 +:temp_w];
assign v496ibus[data_w*2 +:data_w] = c552obus[data_w*1 +:data_w];
assign c552ibus[temp_w*2 +:temp_w] = v730obus[temp_w*2 +:temp_w];
assign v730ibus[data_w*2 +:data_w] = c552obus[data_w*2 +:data_w];
assign c552ibus[temp_w*3 +:temp_w] = v1111obus[temp_w*2 +:temp_w];
assign v1111ibus[data_w*2 +:data_w] = c552obus[data_w*3 +:data_w];
assign c552ibus[temp_w*4 +:temp_w] = v1224obus[temp_w*1 +:temp_w];
assign v1224ibus[data_w*1 +:data_w] = c552obus[data_w*4 +:data_w];
assign c552ibus[temp_w*5 +:temp_w] = v1704obus[temp_w*1 +:temp_w];
assign v1704ibus[data_w*1 +:data_w] = c552obus[data_w*5 +:data_w];
assign c552ibus[temp_w*6 +:temp_w] = v1800obus[temp_w*0 +:temp_w];
assign v1800ibus[data_w*0 +:data_w] = c552obus[data_w*6 +:data_w];
assign c553ibus[temp_w*0 +:temp_w] = v407obus[temp_w*1 +:temp_w];
assign v407ibus[data_w*1 +:data_w] = c553obus[data_w*0 +:data_w];
assign c553ibus[temp_w*1 +:temp_w] = v497obus[temp_w*2 +:temp_w];
assign v497ibus[data_w*2 +:data_w] = c553obus[data_w*1 +:data_w];
assign c553ibus[temp_w*2 +:temp_w] = v731obus[temp_w*2 +:temp_w];
assign v731ibus[data_w*2 +:data_w] = c553obus[data_w*2 +:data_w];
assign c553ibus[temp_w*3 +:temp_w] = v1112obus[temp_w*2 +:temp_w];
assign v1112ibus[data_w*2 +:data_w] = c553obus[data_w*3 +:data_w];
assign c553ibus[temp_w*4 +:temp_w] = v1225obus[temp_w*1 +:temp_w];
assign v1225ibus[data_w*1 +:data_w] = c553obus[data_w*4 +:data_w];
assign c553ibus[temp_w*5 +:temp_w] = v1705obus[temp_w*1 +:temp_w];
assign v1705ibus[data_w*1 +:data_w] = c553obus[data_w*5 +:data_w];
assign c553ibus[temp_w*6 +:temp_w] = v1801obus[temp_w*0 +:temp_w];
assign v1801ibus[data_w*0 +:data_w] = c553obus[data_w*6 +:data_w];
assign c554ibus[temp_w*0 +:temp_w] = v408obus[temp_w*1 +:temp_w];
assign v408ibus[data_w*1 +:data_w] = c554obus[data_w*0 +:data_w];
assign c554ibus[temp_w*1 +:temp_w] = v498obus[temp_w*2 +:temp_w];
assign v498ibus[data_w*2 +:data_w] = c554obus[data_w*1 +:data_w];
assign c554ibus[temp_w*2 +:temp_w] = v732obus[temp_w*2 +:temp_w];
assign v732ibus[data_w*2 +:data_w] = c554obus[data_w*2 +:data_w];
assign c554ibus[temp_w*3 +:temp_w] = v1113obus[temp_w*2 +:temp_w];
assign v1113ibus[data_w*2 +:data_w] = c554obus[data_w*3 +:data_w];
assign c554ibus[temp_w*4 +:temp_w] = v1226obus[temp_w*1 +:temp_w];
assign v1226ibus[data_w*1 +:data_w] = c554obus[data_w*4 +:data_w];
assign c554ibus[temp_w*5 +:temp_w] = v1706obus[temp_w*1 +:temp_w];
assign v1706ibus[data_w*1 +:data_w] = c554obus[data_w*5 +:data_w];
assign c554ibus[temp_w*6 +:temp_w] = v1802obus[temp_w*0 +:temp_w];
assign v1802ibus[data_w*0 +:data_w] = c554obus[data_w*6 +:data_w];
assign c555ibus[temp_w*0 +:temp_w] = v409obus[temp_w*1 +:temp_w];
assign v409ibus[data_w*1 +:data_w] = c555obus[data_w*0 +:data_w];
assign c555ibus[temp_w*1 +:temp_w] = v499obus[temp_w*2 +:temp_w];
assign v499ibus[data_w*2 +:data_w] = c555obus[data_w*1 +:data_w];
assign c555ibus[temp_w*2 +:temp_w] = v733obus[temp_w*2 +:temp_w];
assign v733ibus[data_w*2 +:data_w] = c555obus[data_w*2 +:data_w];
assign c555ibus[temp_w*3 +:temp_w] = v1114obus[temp_w*2 +:temp_w];
assign v1114ibus[data_w*2 +:data_w] = c555obus[data_w*3 +:data_w];
assign c555ibus[temp_w*4 +:temp_w] = v1227obus[temp_w*1 +:temp_w];
assign v1227ibus[data_w*1 +:data_w] = c555obus[data_w*4 +:data_w];
assign c555ibus[temp_w*5 +:temp_w] = v1707obus[temp_w*1 +:temp_w];
assign v1707ibus[data_w*1 +:data_w] = c555obus[data_w*5 +:data_w];
assign c555ibus[temp_w*6 +:temp_w] = v1803obus[temp_w*0 +:temp_w];
assign v1803ibus[data_w*0 +:data_w] = c555obus[data_w*6 +:data_w];
assign c556ibus[temp_w*0 +:temp_w] = v410obus[temp_w*1 +:temp_w];
assign v410ibus[data_w*1 +:data_w] = c556obus[data_w*0 +:data_w];
assign c556ibus[temp_w*1 +:temp_w] = v500obus[temp_w*2 +:temp_w];
assign v500ibus[data_w*2 +:data_w] = c556obus[data_w*1 +:data_w];
assign c556ibus[temp_w*2 +:temp_w] = v734obus[temp_w*2 +:temp_w];
assign v734ibus[data_w*2 +:data_w] = c556obus[data_w*2 +:data_w];
assign c556ibus[temp_w*3 +:temp_w] = v1115obus[temp_w*2 +:temp_w];
assign v1115ibus[data_w*2 +:data_w] = c556obus[data_w*3 +:data_w];
assign c556ibus[temp_w*4 +:temp_w] = v1228obus[temp_w*1 +:temp_w];
assign v1228ibus[data_w*1 +:data_w] = c556obus[data_w*4 +:data_w];
assign c556ibus[temp_w*5 +:temp_w] = v1708obus[temp_w*1 +:temp_w];
assign v1708ibus[data_w*1 +:data_w] = c556obus[data_w*5 +:data_w];
assign c556ibus[temp_w*6 +:temp_w] = v1804obus[temp_w*0 +:temp_w];
assign v1804ibus[data_w*0 +:data_w] = c556obus[data_w*6 +:data_w];
assign c557ibus[temp_w*0 +:temp_w] = v411obus[temp_w*1 +:temp_w];
assign v411ibus[data_w*1 +:data_w] = c557obus[data_w*0 +:data_w];
assign c557ibus[temp_w*1 +:temp_w] = v501obus[temp_w*2 +:temp_w];
assign v501ibus[data_w*2 +:data_w] = c557obus[data_w*1 +:data_w];
assign c557ibus[temp_w*2 +:temp_w] = v735obus[temp_w*2 +:temp_w];
assign v735ibus[data_w*2 +:data_w] = c557obus[data_w*2 +:data_w];
assign c557ibus[temp_w*3 +:temp_w] = v1116obus[temp_w*2 +:temp_w];
assign v1116ibus[data_w*2 +:data_w] = c557obus[data_w*3 +:data_w];
assign c557ibus[temp_w*4 +:temp_w] = v1229obus[temp_w*1 +:temp_w];
assign v1229ibus[data_w*1 +:data_w] = c557obus[data_w*4 +:data_w];
assign c557ibus[temp_w*5 +:temp_w] = v1709obus[temp_w*1 +:temp_w];
assign v1709ibus[data_w*1 +:data_w] = c557obus[data_w*5 +:data_w];
assign c557ibus[temp_w*6 +:temp_w] = v1805obus[temp_w*0 +:temp_w];
assign v1805ibus[data_w*0 +:data_w] = c557obus[data_w*6 +:data_w];
assign c558ibus[temp_w*0 +:temp_w] = v412obus[temp_w*1 +:temp_w];
assign v412ibus[data_w*1 +:data_w] = c558obus[data_w*0 +:data_w];
assign c558ibus[temp_w*1 +:temp_w] = v502obus[temp_w*2 +:temp_w];
assign v502ibus[data_w*2 +:data_w] = c558obus[data_w*1 +:data_w];
assign c558ibus[temp_w*2 +:temp_w] = v736obus[temp_w*2 +:temp_w];
assign v736ibus[data_w*2 +:data_w] = c558obus[data_w*2 +:data_w];
assign c558ibus[temp_w*3 +:temp_w] = v1117obus[temp_w*2 +:temp_w];
assign v1117ibus[data_w*2 +:data_w] = c558obus[data_w*3 +:data_w];
assign c558ibus[temp_w*4 +:temp_w] = v1230obus[temp_w*1 +:temp_w];
assign v1230ibus[data_w*1 +:data_w] = c558obus[data_w*4 +:data_w];
assign c558ibus[temp_w*5 +:temp_w] = v1710obus[temp_w*1 +:temp_w];
assign v1710ibus[data_w*1 +:data_w] = c558obus[data_w*5 +:data_w];
assign c558ibus[temp_w*6 +:temp_w] = v1806obus[temp_w*0 +:temp_w];
assign v1806ibus[data_w*0 +:data_w] = c558obus[data_w*6 +:data_w];
assign c559ibus[temp_w*0 +:temp_w] = v413obus[temp_w*1 +:temp_w];
assign v413ibus[data_w*1 +:data_w] = c559obus[data_w*0 +:data_w];
assign c559ibus[temp_w*1 +:temp_w] = v503obus[temp_w*2 +:temp_w];
assign v503ibus[data_w*2 +:data_w] = c559obus[data_w*1 +:data_w];
assign c559ibus[temp_w*2 +:temp_w] = v737obus[temp_w*2 +:temp_w];
assign v737ibus[data_w*2 +:data_w] = c559obus[data_w*2 +:data_w];
assign c559ibus[temp_w*3 +:temp_w] = v1118obus[temp_w*2 +:temp_w];
assign v1118ibus[data_w*2 +:data_w] = c559obus[data_w*3 +:data_w];
assign c559ibus[temp_w*4 +:temp_w] = v1231obus[temp_w*1 +:temp_w];
assign v1231ibus[data_w*1 +:data_w] = c559obus[data_w*4 +:data_w];
assign c559ibus[temp_w*5 +:temp_w] = v1711obus[temp_w*1 +:temp_w];
assign v1711ibus[data_w*1 +:data_w] = c559obus[data_w*5 +:data_w];
assign c559ibus[temp_w*6 +:temp_w] = v1807obus[temp_w*0 +:temp_w];
assign v1807ibus[data_w*0 +:data_w] = c559obus[data_w*6 +:data_w];
assign c560ibus[temp_w*0 +:temp_w] = v414obus[temp_w*1 +:temp_w];
assign v414ibus[data_w*1 +:data_w] = c560obus[data_w*0 +:data_w];
assign c560ibus[temp_w*1 +:temp_w] = v504obus[temp_w*2 +:temp_w];
assign v504ibus[data_w*2 +:data_w] = c560obus[data_w*1 +:data_w];
assign c560ibus[temp_w*2 +:temp_w] = v738obus[temp_w*2 +:temp_w];
assign v738ibus[data_w*2 +:data_w] = c560obus[data_w*2 +:data_w];
assign c560ibus[temp_w*3 +:temp_w] = v1119obus[temp_w*2 +:temp_w];
assign v1119ibus[data_w*2 +:data_w] = c560obus[data_w*3 +:data_w];
assign c560ibus[temp_w*4 +:temp_w] = v1232obus[temp_w*1 +:temp_w];
assign v1232ibus[data_w*1 +:data_w] = c560obus[data_w*4 +:data_w];
assign c560ibus[temp_w*5 +:temp_w] = v1712obus[temp_w*1 +:temp_w];
assign v1712ibus[data_w*1 +:data_w] = c560obus[data_w*5 +:data_w];
assign c560ibus[temp_w*6 +:temp_w] = v1808obus[temp_w*0 +:temp_w];
assign v1808ibus[data_w*0 +:data_w] = c560obus[data_w*6 +:data_w];
assign c561ibus[temp_w*0 +:temp_w] = v415obus[temp_w*1 +:temp_w];
assign v415ibus[data_w*1 +:data_w] = c561obus[data_w*0 +:data_w];
assign c561ibus[temp_w*1 +:temp_w] = v505obus[temp_w*2 +:temp_w];
assign v505ibus[data_w*2 +:data_w] = c561obus[data_w*1 +:data_w];
assign c561ibus[temp_w*2 +:temp_w] = v739obus[temp_w*2 +:temp_w];
assign v739ibus[data_w*2 +:data_w] = c561obus[data_w*2 +:data_w];
assign c561ibus[temp_w*3 +:temp_w] = v1120obus[temp_w*2 +:temp_w];
assign v1120ibus[data_w*2 +:data_w] = c561obus[data_w*3 +:data_w];
assign c561ibus[temp_w*4 +:temp_w] = v1233obus[temp_w*1 +:temp_w];
assign v1233ibus[data_w*1 +:data_w] = c561obus[data_w*4 +:data_w];
assign c561ibus[temp_w*5 +:temp_w] = v1713obus[temp_w*1 +:temp_w];
assign v1713ibus[data_w*1 +:data_w] = c561obus[data_w*5 +:data_w];
assign c561ibus[temp_w*6 +:temp_w] = v1809obus[temp_w*0 +:temp_w];
assign v1809ibus[data_w*0 +:data_w] = c561obus[data_w*6 +:data_w];
assign c562ibus[temp_w*0 +:temp_w] = v416obus[temp_w*1 +:temp_w];
assign v416ibus[data_w*1 +:data_w] = c562obus[data_w*0 +:data_w];
assign c562ibus[temp_w*1 +:temp_w] = v506obus[temp_w*2 +:temp_w];
assign v506ibus[data_w*2 +:data_w] = c562obus[data_w*1 +:data_w];
assign c562ibus[temp_w*2 +:temp_w] = v740obus[temp_w*2 +:temp_w];
assign v740ibus[data_w*2 +:data_w] = c562obus[data_w*2 +:data_w];
assign c562ibus[temp_w*3 +:temp_w] = v1121obus[temp_w*2 +:temp_w];
assign v1121ibus[data_w*2 +:data_w] = c562obus[data_w*3 +:data_w];
assign c562ibus[temp_w*4 +:temp_w] = v1234obus[temp_w*1 +:temp_w];
assign v1234ibus[data_w*1 +:data_w] = c562obus[data_w*4 +:data_w];
assign c562ibus[temp_w*5 +:temp_w] = v1714obus[temp_w*1 +:temp_w];
assign v1714ibus[data_w*1 +:data_w] = c562obus[data_w*5 +:data_w];
assign c562ibus[temp_w*6 +:temp_w] = v1810obus[temp_w*0 +:temp_w];
assign v1810ibus[data_w*0 +:data_w] = c562obus[data_w*6 +:data_w];
assign c563ibus[temp_w*0 +:temp_w] = v417obus[temp_w*1 +:temp_w];
assign v417ibus[data_w*1 +:data_w] = c563obus[data_w*0 +:data_w];
assign c563ibus[temp_w*1 +:temp_w] = v507obus[temp_w*2 +:temp_w];
assign v507ibus[data_w*2 +:data_w] = c563obus[data_w*1 +:data_w];
assign c563ibus[temp_w*2 +:temp_w] = v741obus[temp_w*2 +:temp_w];
assign v741ibus[data_w*2 +:data_w] = c563obus[data_w*2 +:data_w];
assign c563ibus[temp_w*3 +:temp_w] = v1122obus[temp_w*2 +:temp_w];
assign v1122ibus[data_w*2 +:data_w] = c563obus[data_w*3 +:data_w];
assign c563ibus[temp_w*4 +:temp_w] = v1235obus[temp_w*1 +:temp_w];
assign v1235ibus[data_w*1 +:data_w] = c563obus[data_w*4 +:data_w];
assign c563ibus[temp_w*5 +:temp_w] = v1715obus[temp_w*1 +:temp_w];
assign v1715ibus[data_w*1 +:data_w] = c563obus[data_w*5 +:data_w];
assign c563ibus[temp_w*6 +:temp_w] = v1811obus[temp_w*0 +:temp_w];
assign v1811ibus[data_w*0 +:data_w] = c563obus[data_w*6 +:data_w];
assign c564ibus[temp_w*0 +:temp_w] = v418obus[temp_w*1 +:temp_w];
assign v418ibus[data_w*1 +:data_w] = c564obus[data_w*0 +:data_w];
assign c564ibus[temp_w*1 +:temp_w] = v508obus[temp_w*2 +:temp_w];
assign v508ibus[data_w*2 +:data_w] = c564obus[data_w*1 +:data_w];
assign c564ibus[temp_w*2 +:temp_w] = v742obus[temp_w*2 +:temp_w];
assign v742ibus[data_w*2 +:data_w] = c564obus[data_w*2 +:data_w];
assign c564ibus[temp_w*3 +:temp_w] = v1123obus[temp_w*2 +:temp_w];
assign v1123ibus[data_w*2 +:data_w] = c564obus[data_w*3 +:data_w];
assign c564ibus[temp_w*4 +:temp_w] = v1236obus[temp_w*1 +:temp_w];
assign v1236ibus[data_w*1 +:data_w] = c564obus[data_w*4 +:data_w];
assign c564ibus[temp_w*5 +:temp_w] = v1716obus[temp_w*1 +:temp_w];
assign v1716ibus[data_w*1 +:data_w] = c564obus[data_w*5 +:data_w];
assign c564ibus[temp_w*6 +:temp_w] = v1812obus[temp_w*0 +:temp_w];
assign v1812ibus[data_w*0 +:data_w] = c564obus[data_w*6 +:data_w];
assign c565ibus[temp_w*0 +:temp_w] = v419obus[temp_w*1 +:temp_w];
assign v419ibus[data_w*1 +:data_w] = c565obus[data_w*0 +:data_w];
assign c565ibus[temp_w*1 +:temp_w] = v509obus[temp_w*2 +:temp_w];
assign v509ibus[data_w*2 +:data_w] = c565obus[data_w*1 +:data_w];
assign c565ibus[temp_w*2 +:temp_w] = v743obus[temp_w*2 +:temp_w];
assign v743ibus[data_w*2 +:data_w] = c565obus[data_w*2 +:data_w];
assign c565ibus[temp_w*3 +:temp_w] = v1124obus[temp_w*2 +:temp_w];
assign v1124ibus[data_w*2 +:data_w] = c565obus[data_w*3 +:data_w];
assign c565ibus[temp_w*4 +:temp_w] = v1237obus[temp_w*1 +:temp_w];
assign v1237ibus[data_w*1 +:data_w] = c565obus[data_w*4 +:data_w];
assign c565ibus[temp_w*5 +:temp_w] = v1717obus[temp_w*1 +:temp_w];
assign v1717ibus[data_w*1 +:data_w] = c565obus[data_w*5 +:data_w];
assign c565ibus[temp_w*6 +:temp_w] = v1813obus[temp_w*0 +:temp_w];
assign v1813ibus[data_w*0 +:data_w] = c565obus[data_w*6 +:data_w];
assign c566ibus[temp_w*0 +:temp_w] = v420obus[temp_w*1 +:temp_w];
assign v420ibus[data_w*1 +:data_w] = c566obus[data_w*0 +:data_w];
assign c566ibus[temp_w*1 +:temp_w] = v510obus[temp_w*2 +:temp_w];
assign v510ibus[data_w*2 +:data_w] = c566obus[data_w*1 +:data_w];
assign c566ibus[temp_w*2 +:temp_w] = v744obus[temp_w*2 +:temp_w];
assign v744ibus[data_w*2 +:data_w] = c566obus[data_w*2 +:data_w];
assign c566ibus[temp_w*3 +:temp_w] = v1125obus[temp_w*2 +:temp_w];
assign v1125ibus[data_w*2 +:data_w] = c566obus[data_w*3 +:data_w];
assign c566ibus[temp_w*4 +:temp_w] = v1238obus[temp_w*1 +:temp_w];
assign v1238ibus[data_w*1 +:data_w] = c566obus[data_w*4 +:data_w];
assign c566ibus[temp_w*5 +:temp_w] = v1718obus[temp_w*1 +:temp_w];
assign v1718ibus[data_w*1 +:data_w] = c566obus[data_w*5 +:data_w];
assign c566ibus[temp_w*6 +:temp_w] = v1814obus[temp_w*0 +:temp_w];
assign v1814ibus[data_w*0 +:data_w] = c566obus[data_w*6 +:data_w];
assign c567ibus[temp_w*0 +:temp_w] = v421obus[temp_w*1 +:temp_w];
assign v421ibus[data_w*1 +:data_w] = c567obus[data_w*0 +:data_w];
assign c567ibus[temp_w*1 +:temp_w] = v511obus[temp_w*2 +:temp_w];
assign v511ibus[data_w*2 +:data_w] = c567obus[data_w*1 +:data_w];
assign c567ibus[temp_w*2 +:temp_w] = v745obus[temp_w*2 +:temp_w];
assign v745ibus[data_w*2 +:data_w] = c567obus[data_w*2 +:data_w];
assign c567ibus[temp_w*3 +:temp_w] = v1126obus[temp_w*2 +:temp_w];
assign v1126ibus[data_w*2 +:data_w] = c567obus[data_w*3 +:data_w];
assign c567ibus[temp_w*4 +:temp_w] = v1239obus[temp_w*1 +:temp_w];
assign v1239ibus[data_w*1 +:data_w] = c567obus[data_w*4 +:data_w];
assign c567ibus[temp_w*5 +:temp_w] = v1719obus[temp_w*1 +:temp_w];
assign v1719ibus[data_w*1 +:data_w] = c567obus[data_w*5 +:data_w];
assign c567ibus[temp_w*6 +:temp_w] = v1815obus[temp_w*0 +:temp_w];
assign v1815ibus[data_w*0 +:data_w] = c567obus[data_w*6 +:data_w];
assign c568ibus[temp_w*0 +:temp_w] = v422obus[temp_w*1 +:temp_w];
assign v422ibus[data_w*1 +:data_w] = c568obus[data_w*0 +:data_w];
assign c568ibus[temp_w*1 +:temp_w] = v512obus[temp_w*2 +:temp_w];
assign v512ibus[data_w*2 +:data_w] = c568obus[data_w*1 +:data_w];
assign c568ibus[temp_w*2 +:temp_w] = v746obus[temp_w*2 +:temp_w];
assign v746ibus[data_w*2 +:data_w] = c568obus[data_w*2 +:data_w];
assign c568ibus[temp_w*3 +:temp_w] = v1127obus[temp_w*2 +:temp_w];
assign v1127ibus[data_w*2 +:data_w] = c568obus[data_w*3 +:data_w];
assign c568ibus[temp_w*4 +:temp_w] = v1240obus[temp_w*1 +:temp_w];
assign v1240ibus[data_w*1 +:data_w] = c568obus[data_w*4 +:data_w];
assign c568ibus[temp_w*5 +:temp_w] = v1720obus[temp_w*1 +:temp_w];
assign v1720ibus[data_w*1 +:data_w] = c568obus[data_w*5 +:data_w];
assign c568ibus[temp_w*6 +:temp_w] = v1816obus[temp_w*0 +:temp_w];
assign v1816ibus[data_w*0 +:data_w] = c568obus[data_w*6 +:data_w];
assign c569ibus[temp_w*0 +:temp_w] = v423obus[temp_w*1 +:temp_w];
assign v423ibus[data_w*1 +:data_w] = c569obus[data_w*0 +:data_w];
assign c569ibus[temp_w*1 +:temp_w] = v513obus[temp_w*2 +:temp_w];
assign v513ibus[data_w*2 +:data_w] = c569obus[data_w*1 +:data_w];
assign c569ibus[temp_w*2 +:temp_w] = v747obus[temp_w*2 +:temp_w];
assign v747ibus[data_w*2 +:data_w] = c569obus[data_w*2 +:data_w];
assign c569ibus[temp_w*3 +:temp_w] = v1128obus[temp_w*2 +:temp_w];
assign v1128ibus[data_w*2 +:data_w] = c569obus[data_w*3 +:data_w];
assign c569ibus[temp_w*4 +:temp_w] = v1241obus[temp_w*1 +:temp_w];
assign v1241ibus[data_w*1 +:data_w] = c569obus[data_w*4 +:data_w];
assign c569ibus[temp_w*5 +:temp_w] = v1721obus[temp_w*1 +:temp_w];
assign v1721ibus[data_w*1 +:data_w] = c569obus[data_w*5 +:data_w];
assign c569ibus[temp_w*6 +:temp_w] = v1817obus[temp_w*0 +:temp_w];
assign v1817ibus[data_w*0 +:data_w] = c569obus[data_w*6 +:data_w];
assign c570ibus[temp_w*0 +:temp_w] = v424obus[temp_w*1 +:temp_w];
assign v424ibus[data_w*1 +:data_w] = c570obus[data_w*0 +:data_w];
assign c570ibus[temp_w*1 +:temp_w] = v514obus[temp_w*2 +:temp_w];
assign v514ibus[data_w*2 +:data_w] = c570obus[data_w*1 +:data_w];
assign c570ibus[temp_w*2 +:temp_w] = v748obus[temp_w*2 +:temp_w];
assign v748ibus[data_w*2 +:data_w] = c570obus[data_w*2 +:data_w];
assign c570ibus[temp_w*3 +:temp_w] = v1129obus[temp_w*2 +:temp_w];
assign v1129ibus[data_w*2 +:data_w] = c570obus[data_w*3 +:data_w];
assign c570ibus[temp_w*4 +:temp_w] = v1242obus[temp_w*1 +:temp_w];
assign v1242ibus[data_w*1 +:data_w] = c570obus[data_w*4 +:data_w];
assign c570ibus[temp_w*5 +:temp_w] = v1722obus[temp_w*1 +:temp_w];
assign v1722ibus[data_w*1 +:data_w] = c570obus[data_w*5 +:data_w];
assign c570ibus[temp_w*6 +:temp_w] = v1818obus[temp_w*0 +:temp_w];
assign v1818ibus[data_w*0 +:data_w] = c570obus[data_w*6 +:data_w];
assign c571ibus[temp_w*0 +:temp_w] = v425obus[temp_w*1 +:temp_w];
assign v425ibus[data_w*1 +:data_w] = c571obus[data_w*0 +:data_w];
assign c571ibus[temp_w*1 +:temp_w] = v515obus[temp_w*2 +:temp_w];
assign v515ibus[data_w*2 +:data_w] = c571obus[data_w*1 +:data_w];
assign c571ibus[temp_w*2 +:temp_w] = v749obus[temp_w*2 +:temp_w];
assign v749ibus[data_w*2 +:data_w] = c571obus[data_w*2 +:data_w];
assign c571ibus[temp_w*3 +:temp_w] = v1130obus[temp_w*2 +:temp_w];
assign v1130ibus[data_w*2 +:data_w] = c571obus[data_w*3 +:data_w];
assign c571ibus[temp_w*4 +:temp_w] = v1243obus[temp_w*1 +:temp_w];
assign v1243ibus[data_w*1 +:data_w] = c571obus[data_w*4 +:data_w];
assign c571ibus[temp_w*5 +:temp_w] = v1723obus[temp_w*1 +:temp_w];
assign v1723ibus[data_w*1 +:data_w] = c571obus[data_w*5 +:data_w];
assign c571ibus[temp_w*6 +:temp_w] = v1819obus[temp_w*0 +:temp_w];
assign v1819ibus[data_w*0 +:data_w] = c571obus[data_w*6 +:data_w];
assign c572ibus[temp_w*0 +:temp_w] = v426obus[temp_w*1 +:temp_w];
assign v426ibus[data_w*1 +:data_w] = c572obus[data_w*0 +:data_w];
assign c572ibus[temp_w*1 +:temp_w] = v516obus[temp_w*2 +:temp_w];
assign v516ibus[data_w*2 +:data_w] = c572obus[data_w*1 +:data_w];
assign c572ibus[temp_w*2 +:temp_w] = v750obus[temp_w*2 +:temp_w];
assign v750ibus[data_w*2 +:data_w] = c572obus[data_w*2 +:data_w];
assign c572ibus[temp_w*3 +:temp_w] = v1131obus[temp_w*2 +:temp_w];
assign v1131ibus[data_w*2 +:data_w] = c572obus[data_w*3 +:data_w];
assign c572ibus[temp_w*4 +:temp_w] = v1244obus[temp_w*1 +:temp_w];
assign v1244ibus[data_w*1 +:data_w] = c572obus[data_w*4 +:data_w];
assign c572ibus[temp_w*5 +:temp_w] = v1724obus[temp_w*1 +:temp_w];
assign v1724ibus[data_w*1 +:data_w] = c572obus[data_w*5 +:data_w];
assign c572ibus[temp_w*6 +:temp_w] = v1820obus[temp_w*0 +:temp_w];
assign v1820ibus[data_w*0 +:data_w] = c572obus[data_w*6 +:data_w];
assign c573ibus[temp_w*0 +:temp_w] = v427obus[temp_w*1 +:temp_w];
assign v427ibus[data_w*1 +:data_w] = c573obus[data_w*0 +:data_w];
assign c573ibus[temp_w*1 +:temp_w] = v517obus[temp_w*2 +:temp_w];
assign v517ibus[data_w*2 +:data_w] = c573obus[data_w*1 +:data_w];
assign c573ibus[temp_w*2 +:temp_w] = v751obus[temp_w*2 +:temp_w];
assign v751ibus[data_w*2 +:data_w] = c573obus[data_w*2 +:data_w];
assign c573ibus[temp_w*3 +:temp_w] = v1132obus[temp_w*2 +:temp_w];
assign v1132ibus[data_w*2 +:data_w] = c573obus[data_w*3 +:data_w];
assign c573ibus[temp_w*4 +:temp_w] = v1245obus[temp_w*1 +:temp_w];
assign v1245ibus[data_w*1 +:data_w] = c573obus[data_w*4 +:data_w];
assign c573ibus[temp_w*5 +:temp_w] = v1725obus[temp_w*1 +:temp_w];
assign v1725ibus[data_w*1 +:data_w] = c573obus[data_w*5 +:data_w];
assign c573ibus[temp_w*6 +:temp_w] = v1821obus[temp_w*0 +:temp_w];
assign v1821ibus[data_w*0 +:data_w] = c573obus[data_w*6 +:data_w];
assign c574ibus[temp_w*0 +:temp_w] = v428obus[temp_w*1 +:temp_w];
assign v428ibus[data_w*1 +:data_w] = c574obus[data_w*0 +:data_w];
assign c574ibus[temp_w*1 +:temp_w] = v518obus[temp_w*2 +:temp_w];
assign v518ibus[data_w*2 +:data_w] = c574obus[data_w*1 +:data_w];
assign c574ibus[temp_w*2 +:temp_w] = v752obus[temp_w*2 +:temp_w];
assign v752ibus[data_w*2 +:data_w] = c574obus[data_w*2 +:data_w];
assign c574ibus[temp_w*3 +:temp_w] = v1133obus[temp_w*2 +:temp_w];
assign v1133ibus[data_w*2 +:data_w] = c574obus[data_w*3 +:data_w];
assign c574ibus[temp_w*4 +:temp_w] = v1246obus[temp_w*1 +:temp_w];
assign v1246ibus[data_w*1 +:data_w] = c574obus[data_w*4 +:data_w];
assign c574ibus[temp_w*5 +:temp_w] = v1726obus[temp_w*1 +:temp_w];
assign v1726ibus[data_w*1 +:data_w] = c574obus[data_w*5 +:data_w];
assign c574ibus[temp_w*6 +:temp_w] = v1822obus[temp_w*0 +:temp_w];
assign v1822ibus[data_w*0 +:data_w] = c574obus[data_w*6 +:data_w];
assign c575ibus[temp_w*0 +:temp_w] = v429obus[temp_w*1 +:temp_w];
assign v429ibus[data_w*1 +:data_w] = c575obus[data_w*0 +:data_w];
assign c575ibus[temp_w*1 +:temp_w] = v519obus[temp_w*2 +:temp_w];
assign v519ibus[data_w*2 +:data_w] = c575obus[data_w*1 +:data_w];
assign c575ibus[temp_w*2 +:temp_w] = v753obus[temp_w*2 +:temp_w];
assign v753ibus[data_w*2 +:data_w] = c575obus[data_w*2 +:data_w];
assign c575ibus[temp_w*3 +:temp_w] = v1134obus[temp_w*2 +:temp_w];
assign v1134ibus[data_w*2 +:data_w] = c575obus[data_w*3 +:data_w];
assign c575ibus[temp_w*4 +:temp_w] = v1247obus[temp_w*1 +:temp_w];
assign v1247ibus[data_w*1 +:data_w] = c575obus[data_w*4 +:data_w];
assign c575ibus[temp_w*5 +:temp_w] = v1727obus[temp_w*1 +:temp_w];
assign v1727ibus[data_w*1 +:data_w] = c575obus[data_w*5 +:data_w];
assign c575ibus[temp_w*6 +:temp_w] = v1823obus[temp_w*0 +:temp_w];
assign v1823ibus[data_w*0 +:data_w] = c575obus[data_w*6 +:data_w];
assign c576ibus[temp_w*0 +:temp_w] = v287obus[temp_w*3 +:temp_w];
assign v287ibus[data_w*3 +:data_w] = c576obus[data_w*0 +:data_w];
assign c576ibus[temp_w*1 +:temp_w] = v341obus[temp_w*1 +:temp_w];
assign v341ibus[data_w*1 +:data_w] = c576obus[data_w*1 +:data_w];
assign c576ibus[temp_w*2 +:temp_w] = v878obus[temp_w*3 +:temp_w];
assign v878ibus[data_w*3 +:data_w] = c576obus[data_w*2 +:data_w];
assign c576ibus[temp_w*3 +:temp_w] = v978obus[temp_w*1 +:temp_w];
assign v978ibus[data_w*1 +:data_w] = c576obus[data_w*3 +:data_w];
assign c576ibus[temp_w*4 +:temp_w] = v1728obus[temp_w*1 +:temp_w];
assign v1728ibus[data_w*1 +:data_w] = c576obus[data_w*4 +:data_w];
assign c576ibus[temp_w*5 +:temp_w] = v1824obus[temp_w*0 +:temp_w];
assign v1824ibus[data_w*0 +:data_w] = c576obus[data_w*5 +:data_w];
assign c577ibus[temp_w*0 +:temp_w] = v192obus[temp_w*3 +:temp_w];
assign v192ibus[data_w*3 +:data_w] = c577obus[data_w*0 +:data_w];
assign c577ibus[temp_w*1 +:temp_w] = v342obus[temp_w*1 +:temp_w];
assign v342ibus[data_w*1 +:data_w] = c577obus[data_w*1 +:data_w];
assign c577ibus[temp_w*2 +:temp_w] = v879obus[temp_w*3 +:temp_w];
assign v879ibus[data_w*3 +:data_w] = c577obus[data_w*2 +:data_w];
assign c577ibus[temp_w*3 +:temp_w] = v979obus[temp_w*1 +:temp_w];
assign v979ibus[data_w*1 +:data_w] = c577obus[data_w*3 +:data_w];
assign c577ibus[temp_w*4 +:temp_w] = v1729obus[temp_w*1 +:temp_w];
assign v1729ibus[data_w*1 +:data_w] = c577obus[data_w*4 +:data_w];
assign c577ibus[temp_w*5 +:temp_w] = v1825obus[temp_w*0 +:temp_w];
assign v1825ibus[data_w*0 +:data_w] = c577obus[data_w*5 +:data_w];
assign c578ibus[temp_w*0 +:temp_w] = v193obus[temp_w*3 +:temp_w];
assign v193ibus[data_w*3 +:data_w] = c578obus[data_w*0 +:data_w];
assign c578ibus[temp_w*1 +:temp_w] = v343obus[temp_w*1 +:temp_w];
assign v343ibus[data_w*1 +:data_w] = c578obus[data_w*1 +:data_w];
assign c578ibus[temp_w*2 +:temp_w] = v880obus[temp_w*3 +:temp_w];
assign v880ibus[data_w*3 +:data_w] = c578obus[data_w*2 +:data_w];
assign c578ibus[temp_w*3 +:temp_w] = v980obus[temp_w*1 +:temp_w];
assign v980ibus[data_w*1 +:data_w] = c578obus[data_w*3 +:data_w];
assign c578ibus[temp_w*4 +:temp_w] = v1730obus[temp_w*1 +:temp_w];
assign v1730ibus[data_w*1 +:data_w] = c578obus[data_w*4 +:data_w];
assign c578ibus[temp_w*5 +:temp_w] = v1826obus[temp_w*0 +:temp_w];
assign v1826ibus[data_w*0 +:data_w] = c578obus[data_w*5 +:data_w];
assign c579ibus[temp_w*0 +:temp_w] = v194obus[temp_w*3 +:temp_w];
assign v194ibus[data_w*3 +:data_w] = c579obus[data_w*0 +:data_w];
assign c579ibus[temp_w*1 +:temp_w] = v344obus[temp_w*1 +:temp_w];
assign v344ibus[data_w*1 +:data_w] = c579obus[data_w*1 +:data_w];
assign c579ibus[temp_w*2 +:temp_w] = v881obus[temp_w*3 +:temp_w];
assign v881ibus[data_w*3 +:data_w] = c579obus[data_w*2 +:data_w];
assign c579ibus[temp_w*3 +:temp_w] = v981obus[temp_w*1 +:temp_w];
assign v981ibus[data_w*1 +:data_w] = c579obus[data_w*3 +:data_w];
assign c579ibus[temp_w*4 +:temp_w] = v1731obus[temp_w*1 +:temp_w];
assign v1731ibus[data_w*1 +:data_w] = c579obus[data_w*4 +:data_w];
assign c579ibus[temp_w*5 +:temp_w] = v1827obus[temp_w*0 +:temp_w];
assign v1827ibus[data_w*0 +:data_w] = c579obus[data_w*5 +:data_w];
assign c580ibus[temp_w*0 +:temp_w] = v195obus[temp_w*3 +:temp_w];
assign v195ibus[data_w*3 +:data_w] = c580obus[data_w*0 +:data_w];
assign c580ibus[temp_w*1 +:temp_w] = v345obus[temp_w*1 +:temp_w];
assign v345ibus[data_w*1 +:data_w] = c580obus[data_w*1 +:data_w];
assign c580ibus[temp_w*2 +:temp_w] = v882obus[temp_w*3 +:temp_w];
assign v882ibus[data_w*3 +:data_w] = c580obus[data_w*2 +:data_w];
assign c580ibus[temp_w*3 +:temp_w] = v982obus[temp_w*1 +:temp_w];
assign v982ibus[data_w*1 +:data_w] = c580obus[data_w*3 +:data_w];
assign c580ibus[temp_w*4 +:temp_w] = v1732obus[temp_w*1 +:temp_w];
assign v1732ibus[data_w*1 +:data_w] = c580obus[data_w*4 +:data_w];
assign c580ibus[temp_w*5 +:temp_w] = v1828obus[temp_w*0 +:temp_w];
assign v1828ibus[data_w*0 +:data_w] = c580obus[data_w*5 +:data_w];
assign c581ibus[temp_w*0 +:temp_w] = v196obus[temp_w*3 +:temp_w];
assign v196ibus[data_w*3 +:data_w] = c581obus[data_w*0 +:data_w];
assign c581ibus[temp_w*1 +:temp_w] = v346obus[temp_w*1 +:temp_w];
assign v346ibus[data_w*1 +:data_w] = c581obus[data_w*1 +:data_w];
assign c581ibus[temp_w*2 +:temp_w] = v883obus[temp_w*3 +:temp_w];
assign v883ibus[data_w*3 +:data_w] = c581obus[data_w*2 +:data_w];
assign c581ibus[temp_w*3 +:temp_w] = v983obus[temp_w*1 +:temp_w];
assign v983ibus[data_w*1 +:data_w] = c581obus[data_w*3 +:data_w];
assign c581ibus[temp_w*4 +:temp_w] = v1733obus[temp_w*1 +:temp_w];
assign v1733ibus[data_w*1 +:data_w] = c581obus[data_w*4 +:data_w];
assign c581ibus[temp_w*5 +:temp_w] = v1829obus[temp_w*0 +:temp_w];
assign v1829ibus[data_w*0 +:data_w] = c581obus[data_w*5 +:data_w];
assign c582ibus[temp_w*0 +:temp_w] = v197obus[temp_w*3 +:temp_w];
assign v197ibus[data_w*3 +:data_w] = c582obus[data_w*0 +:data_w];
assign c582ibus[temp_w*1 +:temp_w] = v347obus[temp_w*1 +:temp_w];
assign v347ibus[data_w*1 +:data_w] = c582obus[data_w*1 +:data_w];
assign c582ibus[temp_w*2 +:temp_w] = v884obus[temp_w*3 +:temp_w];
assign v884ibus[data_w*3 +:data_w] = c582obus[data_w*2 +:data_w];
assign c582ibus[temp_w*3 +:temp_w] = v984obus[temp_w*1 +:temp_w];
assign v984ibus[data_w*1 +:data_w] = c582obus[data_w*3 +:data_w];
assign c582ibus[temp_w*4 +:temp_w] = v1734obus[temp_w*1 +:temp_w];
assign v1734ibus[data_w*1 +:data_w] = c582obus[data_w*4 +:data_w];
assign c582ibus[temp_w*5 +:temp_w] = v1830obus[temp_w*0 +:temp_w];
assign v1830ibus[data_w*0 +:data_w] = c582obus[data_w*5 +:data_w];
assign c583ibus[temp_w*0 +:temp_w] = v198obus[temp_w*3 +:temp_w];
assign v198ibus[data_w*3 +:data_w] = c583obus[data_w*0 +:data_w];
assign c583ibus[temp_w*1 +:temp_w] = v348obus[temp_w*1 +:temp_w];
assign v348ibus[data_w*1 +:data_w] = c583obus[data_w*1 +:data_w];
assign c583ibus[temp_w*2 +:temp_w] = v885obus[temp_w*3 +:temp_w];
assign v885ibus[data_w*3 +:data_w] = c583obus[data_w*2 +:data_w];
assign c583ibus[temp_w*3 +:temp_w] = v985obus[temp_w*1 +:temp_w];
assign v985ibus[data_w*1 +:data_w] = c583obus[data_w*3 +:data_w];
assign c583ibus[temp_w*4 +:temp_w] = v1735obus[temp_w*1 +:temp_w];
assign v1735ibus[data_w*1 +:data_w] = c583obus[data_w*4 +:data_w];
assign c583ibus[temp_w*5 +:temp_w] = v1831obus[temp_w*0 +:temp_w];
assign v1831ibus[data_w*0 +:data_w] = c583obus[data_w*5 +:data_w];
assign c584ibus[temp_w*0 +:temp_w] = v199obus[temp_w*3 +:temp_w];
assign v199ibus[data_w*3 +:data_w] = c584obus[data_w*0 +:data_w];
assign c584ibus[temp_w*1 +:temp_w] = v349obus[temp_w*1 +:temp_w];
assign v349ibus[data_w*1 +:data_w] = c584obus[data_w*1 +:data_w];
assign c584ibus[temp_w*2 +:temp_w] = v886obus[temp_w*3 +:temp_w];
assign v886ibus[data_w*3 +:data_w] = c584obus[data_w*2 +:data_w];
assign c584ibus[temp_w*3 +:temp_w] = v986obus[temp_w*1 +:temp_w];
assign v986ibus[data_w*1 +:data_w] = c584obus[data_w*3 +:data_w];
assign c584ibus[temp_w*4 +:temp_w] = v1736obus[temp_w*1 +:temp_w];
assign v1736ibus[data_w*1 +:data_w] = c584obus[data_w*4 +:data_w];
assign c584ibus[temp_w*5 +:temp_w] = v1832obus[temp_w*0 +:temp_w];
assign v1832ibus[data_w*0 +:data_w] = c584obus[data_w*5 +:data_w];
assign c585ibus[temp_w*0 +:temp_w] = v200obus[temp_w*3 +:temp_w];
assign v200ibus[data_w*3 +:data_w] = c585obus[data_w*0 +:data_w];
assign c585ibus[temp_w*1 +:temp_w] = v350obus[temp_w*1 +:temp_w];
assign v350ibus[data_w*1 +:data_w] = c585obus[data_w*1 +:data_w];
assign c585ibus[temp_w*2 +:temp_w] = v887obus[temp_w*3 +:temp_w];
assign v887ibus[data_w*3 +:data_w] = c585obus[data_w*2 +:data_w];
assign c585ibus[temp_w*3 +:temp_w] = v987obus[temp_w*1 +:temp_w];
assign v987ibus[data_w*1 +:data_w] = c585obus[data_w*3 +:data_w];
assign c585ibus[temp_w*4 +:temp_w] = v1737obus[temp_w*1 +:temp_w];
assign v1737ibus[data_w*1 +:data_w] = c585obus[data_w*4 +:data_w];
assign c585ibus[temp_w*5 +:temp_w] = v1833obus[temp_w*0 +:temp_w];
assign v1833ibus[data_w*0 +:data_w] = c585obus[data_w*5 +:data_w];
assign c586ibus[temp_w*0 +:temp_w] = v201obus[temp_w*3 +:temp_w];
assign v201ibus[data_w*3 +:data_w] = c586obus[data_w*0 +:data_w];
assign c586ibus[temp_w*1 +:temp_w] = v351obus[temp_w*1 +:temp_w];
assign v351ibus[data_w*1 +:data_w] = c586obus[data_w*1 +:data_w];
assign c586ibus[temp_w*2 +:temp_w] = v888obus[temp_w*3 +:temp_w];
assign v888ibus[data_w*3 +:data_w] = c586obus[data_w*2 +:data_w];
assign c586ibus[temp_w*3 +:temp_w] = v988obus[temp_w*1 +:temp_w];
assign v988ibus[data_w*1 +:data_w] = c586obus[data_w*3 +:data_w];
assign c586ibus[temp_w*4 +:temp_w] = v1738obus[temp_w*1 +:temp_w];
assign v1738ibus[data_w*1 +:data_w] = c586obus[data_w*4 +:data_w];
assign c586ibus[temp_w*5 +:temp_w] = v1834obus[temp_w*0 +:temp_w];
assign v1834ibus[data_w*0 +:data_w] = c586obus[data_w*5 +:data_w];
assign c587ibus[temp_w*0 +:temp_w] = v202obus[temp_w*3 +:temp_w];
assign v202ibus[data_w*3 +:data_w] = c587obus[data_w*0 +:data_w];
assign c587ibus[temp_w*1 +:temp_w] = v352obus[temp_w*1 +:temp_w];
assign v352ibus[data_w*1 +:data_w] = c587obus[data_w*1 +:data_w];
assign c587ibus[temp_w*2 +:temp_w] = v889obus[temp_w*3 +:temp_w];
assign v889ibus[data_w*3 +:data_w] = c587obus[data_w*2 +:data_w];
assign c587ibus[temp_w*3 +:temp_w] = v989obus[temp_w*1 +:temp_w];
assign v989ibus[data_w*1 +:data_w] = c587obus[data_w*3 +:data_w];
assign c587ibus[temp_w*4 +:temp_w] = v1739obus[temp_w*1 +:temp_w];
assign v1739ibus[data_w*1 +:data_w] = c587obus[data_w*4 +:data_w];
assign c587ibus[temp_w*5 +:temp_w] = v1835obus[temp_w*0 +:temp_w];
assign v1835ibus[data_w*0 +:data_w] = c587obus[data_w*5 +:data_w];
assign c588ibus[temp_w*0 +:temp_w] = v203obus[temp_w*3 +:temp_w];
assign v203ibus[data_w*3 +:data_w] = c588obus[data_w*0 +:data_w];
assign c588ibus[temp_w*1 +:temp_w] = v353obus[temp_w*1 +:temp_w];
assign v353ibus[data_w*1 +:data_w] = c588obus[data_w*1 +:data_w];
assign c588ibus[temp_w*2 +:temp_w] = v890obus[temp_w*3 +:temp_w];
assign v890ibus[data_w*3 +:data_w] = c588obus[data_w*2 +:data_w];
assign c588ibus[temp_w*3 +:temp_w] = v990obus[temp_w*1 +:temp_w];
assign v990ibus[data_w*1 +:data_w] = c588obus[data_w*3 +:data_w];
assign c588ibus[temp_w*4 +:temp_w] = v1740obus[temp_w*1 +:temp_w];
assign v1740ibus[data_w*1 +:data_w] = c588obus[data_w*4 +:data_w];
assign c588ibus[temp_w*5 +:temp_w] = v1836obus[temp_w*0 +:temp_w];
assign v1836ibus[data_w*0 +:data_w] = c588obus[data_w*5 +:data_w];
assign c589ibus[temp_w*0 +:temp_w] = v204obus[temp_w*3 +:temp_w];
assign v204ibus[data_w*3 +:data_w] = c589obus[data_w*0 +:data_w];
assign c589ibus[temp_w*1 +:temp_w] = v354obus[temp_w*1 +:temp_w];
assign v354ibus[data_w*1 +:data_w] = c589obus[data_w*1 +:data_w];
assign c589ibus[temp_w*2 +:temp_w] = v891obus[temp_w*3 +:temp_w];
assign v891ibus[data_w*3 +:data_w] = c589obus[data_w*2 +:data_w];
assign c589ibus[temp_w*3 +:temp_w] = v991obus[temp_w*1 +:temp_w];
assign v991ibus[data_w*1 +:data_w] = c589obus[data_w*3 +:data_w];
assign c589ibus[temp_w*4 +:temp_w] = v1741obus[temp_w*1 +:temp_w];
assign v1741ibus[data_w*1 +:data_w] = c589obus[data_w*4 +:data_w];
assign c589ibus[temp_w*5 +:temp_w] = v1837obus[temp_w*0 +:temp_w];
assign v1837ibus[data_w*0 +:data_w] = c589obus[data_w*5 +:data_w];
assign c590ibus[temp_w*0 +:temp_w] = v205obus[temp_w*3 +:temp_w];
assign v205ibus[data_w*3 +:data_w] = c590obus[data_w*0 +:data_w];
assign c590ibus[temp_w*1 +:temp_w] = v355obus[temp_w*1 +:temp_w];
assign v355ibus[data_w*1 +:data_w] = c590obus[data_w*1 +:data_w];
assign c590ibus[temp_w*2 +:temp_w] = v892obus[temp_w*3 +:temp_w];
assign v892ibus[data_w*3 +:data_w] = c590obus[data_w*2 +:data_w];
assign c590ibus[temp_w*3 +:temp_w] = v992obus[temp_w*1 +:temp_w];
assign v992ibus[data_w*1 +:data_w] = c590obus[data_w*3 +:data_w];
assign c590ibus[temp_w*4 +:temp_w] = v1742obus[temp_w*1 +:temp_w];
assign v1742ibus[data_w*1 +:data_w] = c590obus[data_w*4 +:data_w];
assign c590ibus[temp_w*5 +:temp_w] = v1838obus[temp_w*0 +:temp_w];
assign v1838ibus[data_w*0 +:data_w] = c590obus[data_w*5 +:data_w];
assign c591ibus[temp_w*0 +:temp_w] = v206obus[temp_w*3 +:temp_w];
assign v206ibus[data_w*3 +:data_w] = c591obus[data_w*0 +:data_w];
assign c591ibus[temp_w*1 +:temp_w] = v356obus[temp_w*1 +:temp_w];
assign v356ibus[data_w*1 +:data_w] = c591obus[data_w*1 +:data_w];
assign c591ibus[temp_w*2 +:temp_w] = v893obus[temp_w*3 +:temp_w];
assign v893ibus[data_w*3 +:data_w] = c591obus[data_w*2 +:data_w];
assign c591ibus[temp_w*3 +:temp_w] = v993obus[temp_w*1 +:temp_w];
assign v993ibus[data_w*1 +:data_w] = c591obus[data_w*3 +:data_w];
assign c591ibus[temp_w*4 +:temp_w] = v1743obus[temp_w*1 +:temp_w];
assign v1743ibus[data_w*1 +:data_w] = c591obus[data_w*4 +:data_w];
assign c591ibus[temp_w*5 +:temp_w] = v1839obus[temp_w*0 +:temp_w];
assign v1839ibus[data_w*0 +:data_w] = c591obus[data_w*5 +:data_w];
assign c592ibus[temp_w*0 +:temp_w] = v207obus[temp_w*3 +:temp_w];
assign v207ibus[data_w*3 +:data_w] = c592obus[data_w*0 +:data_w];
assign c592ibus[temp_w*1 +:temp_w] = v357obus[temp_w*1 +:temp_w];
assign v357ibus[data_w*1 +:data_w] = c592obus[data_w*1 +:data_w];
assign c592ibus[temp_w*2 +:temp_w] = v894obus[temp_w*3 +:temp_w];
assign v894ibus[data_w*3 +:data_w] = c592obus[data_w*2 +:data_w];
assign c592ibus[temp_w*3 +:temp_w] = v994obus[temp_w*1 +:temp_w];
assign v994ibus[data_w*1 +:data_w] = c592obus[data_w*3 +:data_w];
assign c592ibus[temp_w*4 +:temp_w] = v1744obus[temp_w*1 +:temp_w];
assign v1744ibus[data_w*1 +:data_w] = c592obus[data_w*4 +:data_w];
assign c592ibus[temp_w*5 +:temp_w] = v1840obus[temp_w*0 +:temp_w];
assign v1840ibus[data_w*0 +:data_w] = c592obus[data_w*5 +:data_w];
assign c593ibus[temp_w*0 +:temp_w] = v208obus[temp_w*3 +:temp_w];
assign v208ibus[data_w*3 +:data_w] = c593obus[data_w*0 +:data_w];
assign c593ibus[temp_w*1 +:temp_w] = v358obus[temp_w*1 +:temp_w];
assign v358ibus[data_w*1 +:data_w] = c593obus[data_w*1 +:data_w];
assign c593ibus[temp_w*2 +:temp_w] = v895obus[temp_w*3 +:temp_w];
assign v895ibus[data_w*3 +:data_w] = c593obus[data_w*2 +:data_w];
assign c593ibus[temp_w*3 +:temp_w] = v995obus[temp_w*1 +:temp_w];
assign v995ibus[data_w*1 +:data_w] = c593obus[data_w*3 +:data_w];
assign c593ibus[temp_w*4 +:temp_w] = v1745obus[temp_w*1 +:temp_w];
assign v1745ibus[data_w*1 +:data_w] = c593obus[data_w*4 +:data_w];
assign c593ibus[temp_w*5 +:temp_w] = v1841obus[temp_w*0 +:temp_w];
assign v1841ibus[data_w*0 +:data_w] = c593obus[data_w*5 +:data_w];
assign c594ibus[temp_w*0 +:temp_w] = v209obus[temp_w*3 +:temp_w];
assign v209ibus[data_w*3 +:data_w] = c594obus[data_w*0 +:data_w];
assign c594ibus[temp_w*1 +:temp_w] = v359obus[temp_w*1 +:temp_w];
assign v359ibus[data_w*1 +:data_w] = c594obus[data_w*1 +:data_w];
assign c594ibus[temp_w*2 +:temp_w] = v896obus[temp_w*3 +:temp_w];
assign v896ibus[data_w*3 +:data_w] = c594obus[data_w*2 +:data_w];
assign c594ibus[temp_w*3 +:temp_w] = v996obus[temp_w*1 +:temp_w];
assign v996ibus[data_w*1 +:data_w] = c594obus[data_w*3 +:data_w];
assign c594ibus[temp_w*4 +:temp_w] = v1746obus[temp_w*1 +:temp_w];
assign v1746ibus[data_w*1 +:data_w] = c594obus[data_w*4 +:data_w];
assign c594ibus[temp_w*5 +:temp_w] = v1842obus[temp_w*0 +:temp_w];
assign v1842ibus[data_w*0 +:data_w] = c594obus[data_w*5 +:data_w];
assign c595ibus[temp_w*0 +:temp_w] = v210obus[temp_w*3 +:temp_w];
assign v210ibus[data_w*3 +:data_w] = c595obus[data_w*0 +:data_w];
assign c595ibus[temp_w*1 +:temp_w] = v360obus[temp_w*1 +:temp_w];
assign v360ibus[data_w*1 +:data_w] = c595obus[data_w*1 +:data_w];
assign c595ibus[temp_w*2 +:temp_w] = v897obus[temp_w*3 +:temp_w];
assign v897ibus[data_w*3 +:data_w] = c595obus[data_w*2 +:data_w];
assign c595ibus[temp_w*3 +:temp_w] = v997obus[temp_w*1 +:temp_w];
assign v997ibus[data_w*1 +:data_w] = c595obus[data_w*3 +:data_w];
assign c595ibus[temp_w*4 +:temp_w] = v1747obus[temp_w*1 +:temp_w];
assign v1747ibus[data_w*1 +:data_w] = c595obus[data_w*4 +:data_w];
assign c595ibus[temp_w*5 +:temp_w] = v1843obus[temp_w*0 +:temp_w];
assign v1843ibus[data_w*0 +:data_w] = c595obus[data_w*5 +:data_w];
assign c596ibus[temp_w*0 +:temp_w] = v211obus[temp_w*3 +:temp_w];
assign v211ibus[data_w*3 +:data_w] = c596obus[data_w*0 +:data_w];
assign c596ibus[temp_w*1 +:temp_w] = v361obus[temp_w*1 +:temp_w];
assign v361ibus[data_w*1 +:data_w] = c596obus[data_w*1 +:data_w];
assign c596ibus[temp_w*2 +:temp_w] = v898obus[temp_w*3 +:temp_w];
assign v898ibus[data_w*3 +:data_w] = c596obus[data_w*2 +:data_w];
assign c596ibus[temp_w*3 +:temp_w] = v998obus[temp_w*1 +:temp_w];
assign v998ibus[data_w*1 +:data_w] = c596obus[data_w*3 +:data_w];
assign c596ibus[temp_w*4 +:temp_w] = v1748obus[temp_w*1 +:temp_w];
assign v1748ibus[data_w*1 +:data_w] = c596obus[data_w*4 +:data_w];
assign c596ibus[temp_w*5 +:temp_w] = v1844obus[temp_w*0 +:temp_w];
assign v1844ibus[data_w*0 +:data_w] = c596obus[data_w*5 +:data_w];
assign c597ibus[temp_w*0 +:temp_w] = v212obus[temp_w*3 +:temp_w];
assign v212ibus[data_w*3 +:data_w] = c597obus[data_w*0 +:data_w];
assign c597ibus[temp_w*1 +:temp_w] = v362obus[temp_w*1 +:temp_w];
assign v362ibus[data_w*1 +:data_w] = c597obus[data_w*1 +:data_w];
assign c597ibus[temp_w*2 +:temp_w] = v899obus[temp_w*3 +:temp_w];
assign v899ibus[data_w*3 +:data_w] = c597obus[data_w*2 +:data_w];
assign c597ibus[temp_w*3 +:temp_w] = v999obus[temp_w*1 +:temp_w];
assign v999ibus[data_w*1 +:data_w] = c597obus[data_w*3 +:data_w];
assign c597ibus[temp_w*4 +:temp_w] = v1749obus[temp_w*1 +:temp_w];
assign v1749ibus[data_w*1 +:data_w] = c597obus[data_w*4 +:data_w];
assign c597ibus[temp_w*5 +:temp_w] = v1845obus[temp_w*0 +:temp_w];
assign v1845ibus[data_w*0 +:data_w] = c597obus[data_w*5 +:data_w];
assign c598ibus[temp_w*0 +:temp_w] = v213obus[temp_w*3 +:temp_w];
assign v213ibus[data_w*3 +:data_w] = c598obus[data_w*0 +:data_w];
assign c598ibus[temp_w*1 +:temp_w] = v363obus[temp_w*1 +:temp_w];
assign v363ibus[data_w*1 +:data_w] = c598obus[data_w*1 +:data_w];
assign c598ibus[temp_w*2 +:temp_w] = v900obus[temp_w*3 +:temp_w];
assign v900ibus[data_w*3 +:data_w] = c598obus[data_w*2 +:data_w];
assign c598ibus[temp_w*3 +:temp_w] = v1000obus[temp_w*1 +:temp_w];
assign v1000ibus[data_w*1 +:data_w] = c598obus[data_w*3 +:data_w];
assign c598ibus[temp_w*4 +:temp_w] = v1750obus[temp_w*1 +:temp_w];
assign v1750ibus[data_w*1 +:data_w] = c598obus[data_w*4 +:data_w];
assign c598ibus[temp_w*5 +:temp_w] = v1846obus[temp_w*0 +:temp_w];
assign v1846ibus[data_w*0 +:data_w] = c598obus[data_w*5 +:data_w];
assign c599ibus[temp_w*0 +:temp_w] = v214obus[temp_w*3 +:temp_w];
assign v214ibus[data_w*3 +:data_w] = c599obus[data_w*0 +:data_w];
assign c599ibus[temp_w*1 +:temp_w] = v364obus[temp_w*1 +:temp_w];
assign v364ibus[data_w*1 +:data_w] = c599obus[data_w*1 +:data_w];
assign c599ibus[temp_w*2 +:temp_w] = v901obus[temp_w*3 +:temp_w];
assign v901ibus[data_w*3 +:data_w] = c599obus[data_w*2 +:data_w];
assign c599ibus[temp_w*3 +:temp_w] = v1001obus[temp_w*1 +:temp_w];
assign v1001ibus[data_w*1 +:data_w] = c599obus[data_w*3 +:data_w];
assign c599ibus[temp_w*4 +:temp_w] = v1751obus[temp_w*1 +:temp_w];
assign v1751ibus[data_w*1 +:data_w] = c599obus[data_w*4 +:data_w];
assign c599ibus[temp_w*5 +:temp_w] = v1847obus[temp_w*0 +:temp_w];
assign v1847ibus[data_w*0 +:data_w] = c599obus[data_w*5 +:data_w];
assign c600ibus[temp_w*0 +:temp_w] = v215obus[temp_w*3 +:temp_w];
assign v215ibus[data_w*3 +:data_w] = c600obus[data_w*0 +:data_w];
assign c600ibus[temp_w*1 +:temp_w] = v365obus[temp_w*1 +:temp_w];
assign v365ibus[data_w*1 +:data_w] = c600obus[data_w*1 +:data_w];
assign c600ibus[temp_w*2 +:temp_w] = v902obus[temp_w*3 +:temp_w];
assign v902ibus[data_w*3 +:data_w] = c600obus[data_w*2 +:data_w];
assign c600ibus[temp_w*3 +:temp_w] = v1002obus[temp_w*1 +:temp_w];
assign v1002ibus[data_w*1 +:data_w] = c600obus[data_w*3 +:data_w];
assign c600ibus[temp_w*4 +:temp_w] = v1752obus[temp_w*1 +:temp_w];
assign v1752ibus[data_w*1 +:data_w] = c600obus[data_w*4 +:data_w];
assign c600ibus[temp_w*5 +:temp_w] = v1848obus[temp_w*0 +:temp_w];
assign v1848ibus[data_w*0 +:data_w] = c600obus[data_w*5 +:data_w];
assign c601ibus[temp_w*0 +:temp_w] = v216obus[temp_w*3 +:temp_w];
assign v216ibus[data_w*3 +:data_w] = c601obus[data_w*0 +:data_w];
assign c601ibus[temp_w*1 +:temp_w] = v366obus[temp_w*1 +:temp_w];
assign v366ibus[data_w*1 +:data_w] = c601obus[data_w*1 +:data_w];
assign c601ibus[temp_w*2 +:temp_w] = v903obus[temp_w*3 +:temp_w];
assign v903ibus[data_w*3 +:data_w] = c601obus[data_w*2 +:data_w];
assign c601ibus[temp_w*3 +:temp_w] = v1003obus[temp_w*1 +:temp_w];
assign v1003ibus[data_w*1 +:data_w] = c601obus[data_w*3 +:data_w];
assign c601ibus[temp_w*4 +:temp_w] = v1753obus[temp_w*1 +:temp_w];
assign v1753ibus[data_w*1 +:data_w] = c601obus[data_w*4 +:data_w];
assign c601ibus[temp_w*5 +:temp_w] = v1849obus[temp_w*0 +:temp_w];
assign v1849ibus[data_w*0 +:data_w] = c601obus[data_w*5 +:data_w];
assign c602ibus[temp_w*0 +:temp_w] = v217obus[temp_w*3 +:temp_w];
assign v217ibus[data_w*3 +:data_w] = c602obus[data_w*0 +:data_w];
assign c602ibus[temp_w*1 +:temp_w] = v367obus[temp_w*1 +:temp_w];
assign v367ibus[data_w*1 +:data_w] = c602obus[data_w*1 +:data_w];
assign c602ibus[temp_w*2 +:temp_w] = v904obus[temp_w*3 +:temp_w];
assign v904ibus[data_w*3 +:data_w] = c602obus[data_w*2 +:data_w];
assign c602ibus[temp_w*3 +:temp_w] = v1004obus[temp_w*1 +:temp_w];
assign v1004ibus[data_w*1 +:data_w] = c602obus[data_w*3 +:data_w];
assign c602ibus[temp_w*4 +:temp_w] = v1754obus[temp_w*1 +:temp_w];
assign v1754ibus[data_w*1 +:data_w] = c602obus[data_w*4 +:data_w];
assign c602ibus[temp_w*5 +:temp_w] = v1850obus[temp_w*0 +:temp_w];
assign v1850ibus[data_w*0 +:data_w] = c602obus[data_w*5 +:data_w];
assign c603ibus[temp_w*0 +:temp_w] = v218obus[temp_w*3 +:temp_w];
assign v218ibus[data_w*3 +:data_w] = c603obus[data_w*0 +:data_w];
assign c603ibus[temp_w*1 +:temp_w] = v368obus[temp_w*1 +:temp_w];
assign v368ibus[data_w*1 +:data_w] = c603obus[data_w*1 +:data_w];
assign c603ibus[temp_w*2 +:temp_w] = v905obus[temp_w*3 +:temp_w];
assign v905ibus[data_w*3 +:data_w] = c603obus[data_w*2 +:data_w];
assign c603ibus[temp_w*3 +:temp_w] = v1005obus[temp_w*1 +:temp_w];
assign v1005ibus[data_w*1 +:data_w] = c603obus[data_w*3 +:data_w];
assign c603ibus[temp_w*4 +:temp_w] = v1755obus[temp_w*1 +:temp_w];
assign v1755ibus[data_w*1 +:data_w] = c603obus[data_w*4 +:data_w];
assign c603ibus[temp_w*5 +:temp_w] = v1851obus[temp_w*0 +:temp_w];
assign v1851ibus[data_w*0 +:data_w] = c603obus[data_w*5 +:data_w];
assign c604ibus[temp_w*0 +:temp_w] = v219obus[temp_w*3 +:temp_w];
assign v219ibus[data_w*3 +:data_w] = c604obus[data_w*0 +:data_w];
assign c604ibus[temp_w*1 +:temp_w] = v369obus[temp_w*1 +:temp_w];
assign v369ibus[data_w*1 +:data_w] = c604obus[data_w*1 +:data_w];
assign c604ibus[temp_w*2 +:temp_w] = v906obus[temp_w*3 +:temp_w];
assign v906ibus[data_w*3 +:data_w] = c604obus[data_w*2 +:data_w];
assign c604ibus[temp_w*3 +:temp_w] = v1006obus[temp_w*1 +:temp_w];
assign v1006ibus[data_w*1 +:data_w] = c604obus[data_w*3 +:data_w];
assign c604ibus[temp_w*4 +:temp_w] = v1756obus[temp_w*1 +:temp_w];
assign v1756ibus[data_w*1 +:data_w] = c604obus[data_w*4 +:data_w];
assign c604ibus[temp_w*5 +:temp_w] = v1852obus[temp_w*0 +:temp_w];
assign v1852ibus[data_w*0 +:data_w] = c604obus[data_w*5 +:data_w];
assign c605ibus[temp_w*0 +:temp_w] = v220obus[temp_w*3 +:temp_w];
assign v220ibus[data_w*3 +:data_w] = c605obus[data_w*0 +:data_w];
assign c605ibus[temp_w*1 +:temp_w] = v370obus[temp_w*1 +:temp_w];
assign v370ibus[data_w*1 +:data_w] = c605obus[data_w*1 +:data_w];
assign c605ibus[temp_w*2 +:temp_w] = v907obus[temp_w*3 +:temp_w];
assign v907ibus[data_w*3 +:data_w] = c605obus[data_w*2 +:data_w];
assign c605ibus[temp_w*3 +:temp_w] = v1007obus[temp_w*1 +:temp_w];
assign v1007ibus[data_w*1 +:data_w] = c605obus[data_w*3 +:data_w];
assign c605ibus[temp_w*4 +:temp_w] = v1757obus[temp_w*1 +:temp_w];
assign v1757ibus[data_w*1 +:data_w] = c605obus[data_w*4 +:data_w];
assign c605ibus[temp_w*5 +:temp_w] = v1853obus[temp_w*0 +:temp_w];
assign v1853ibus[data_w*0 +:data_w] = c605obus[data_w*5 +:data_w];
assign c606ibus[temp_w*0 +:temp_w] = v221obus[temp_w*3 +:temp_w];
assign v221ibus[data_w*3 +:data_w] = c606obus[data_w*0 +:data_w];
assign c606ibus[temp_w*1 +:temp_w] = v371obus[temp_w*1 +:temp_w];
assign v371ibus[data_w*1 +:data_w] = c606obus[data_w*1 +:data_w];
assign c606ibus[temp_w*2 +:temp_w] = v908obus[temp_w*3 +:temp_w];
assign v908ibus[data_w*3 +:data_w] = c606obus[data_w*2 +:data_w];
assign c606ibus[temp_w*3 +:temp_w] = v1008obus[temp_w*1 +:temp_w];
assign v1008ibus[data_w*1 +:data_w] = c606obus[data_w*3 +:data_w];
assign c606ibus[temp_w*4 +:temp_w] = v1758obus[temp_w*1 +:temp_w];
assign v1758ibus[data_w*1 +:data_w] = c606obus[data_w*4 +:data_w];
assign c606ibus[temp_w*5 +:temp_w] = v1854obus[temp_w*0 +:temp_w];
assign v1854ibus[data_w*0 +:data_w] = c606obus[data_w*5 +:data_w];
assign c607ibus[temp_w*0 +:temp_w] = v222obus[temp_w*3 +:temp_w];
assign v222ibus[data_w*3 +:data_w] = c607obus[data_w*0 +:data_w];
assign c607ibus[temp_w*1 +:temp_w] = v372obus[temp_w*1 +:temp_w];
assign v372ibus[data_w*1 +:data_w] = c607obus[data_w*1 +:data_w];
assign c607ibus[temp_w*2 +:temp_w] = v909obus[temp_w*3 +:temp_w];
assign v909ibus[data_w*3 +:data_w] = c607obus[data_w*2 +:data_w];
assign c607ibus[temp_w*3 +:temp_w] = v1009obus[temp_w*1 +:temp_w];
assign v1009ibus[data_w*1 +:data_w] = c607obus[data_w*3 +:data_w];
assign c607ibus[temp_w*4 +:temp_w] = v1759obus[temp_w*1 +:temp_w];
assign v1759ibus[data_w*1 +:data_w] = c607obus[data_w*4 +:data_w];
assign c607ibus[temp_w*5 +:temp_w] = v1855obus[temp_w*0 +:temp_w];
assign v1855ibus[data_w*0 +:data_w] = c607obus[data_w*5 +:data_w];
assign c608ibus[temp_w*0 +:temp_w] = v223obus[temp_w*3 +:temp_w];
assign v223ibus[data_w*3 +:data_w] = c608obus[data_w*0 +:data_w];
assign c608ibus[temp_w*1 +:temp_w] = v373obus[temp_w*1 +:temp_w];
assign v373ibus[data_w*1 +:data_w] = c608obus[data_w*1 +:data_w];
assign c608ibus[temp_w*2 +:temp_w] = v910obus[temp_w*3 +:temp_w];
assign v910ibus[data_w*3 +:data_w] = c608obus[data_w*2 +:data_w];
assign c608ibus[temp_w*3 +:temp_w] = v1010obus[temp_w*1 +:temp_w];
assign v1010ibus[data_w*1 +:data_w] = c608obus[data_w*3 +:data_w];
assign c608ibus[temp_w*4 +:temp_w] = v1760obus[temp_w*1 +:temp_w];
assign v1760ibus[data_w*1 +:data_w] = c608obus[data_w*4 +:data_w];
assign c608ibus[temp_w*5 +:temp_w] = v1856obus[temp_w*0 +:temp_w];
assign v1856ibus[data_w*0 +:data_w] = c608obus[data_w*5 +:data_w];
assign c609ibus[temp_w*0 +:temp_w] = v224obus[temp_w*3 +:temp_w];
assign v224ibus[data_w*3 +:data_w] = c609obus[data_w*0 +:data_w];
assign c609ibus[temp_w*1 +:temp_w] = v374obus[temp_w*1 +:temp_w];
assign v374ibus[data_w*1 +:data_w] = c609obus[data_w*1 +:data_w];
assign c609ibus[temp_w*2 +:temp_w] = v911obus[temp_w*3 +:temp_w];
assign v911ibus[data_w*3 +:data_w] = c609obus[data_w*2 +:data_w];
assign c609ibus[temp_w*3 +:temp_w] = v1011obus[temp_w*1 +:temp_w];
assign v1011ibus[data_w*1 +:data_w] = c609obus[data_w*3 +:data_w];
assign c609ibus[temp_w*4 +:temp_w] = v1761obus[temp_w*1 +:temp_w];
assign v1761ibus[data_w*1 +:data_w] = c609obus[data_w*4 +:data_w];
assign c609ibus[temp_w*5 +:temp_w] = v1857obus[temp_w*0 +:temp_w];
assign v1857ibus[data_w*0 +:data_w] = c609obus[data_w*5 +:data_w];
assign c610ibus[temp_w*0 +:temp_w] = v225obus[temp_w*3 +:temp_w];
assign v225ibus[data_w*3 +:data_w] = c610obus[data_w*0 +:data_w];
assign c610ibus[temp_w*1 +:temp_w] = v375obus[temp_w*1 +:temp_w];
assign v375ibus[data_w*1 +:data_w] = c610obus[data_w*1 +:data_w];
assign c610ibus[temp_w*2 +:temp_w] = v912obus[temp_w*3 +:temp_w];
assign v912ibus[data_w*3 +:data_w] = c610obus[data_w*2 +:data_w];
assign c610ibus[temp_w*3 +:temp_w] = v1012obus[temp_w*1 +:temp_w];
assign v1012ibus[data_w*1 +:data_w] = c610obus[data_w*3 +:data_w];
assign c610ibus[temp_w*4 +:temp_w] = v1762obus[temp_w*1 +:temp_w];
assign v1762ibus[data_w*1 +:data_w] = c610obus[data_w*4 +:data_w];
assign c610ibus[temp_w*5 +:temp_w] = v1858obus[temp_w*0 +:temp_w];
assign v1858ibus[data_w*0 +:data_w] = c610obus[data_w*5 +:data_w];
assign c611ibus[temp_w*0 +:temp_w] = v226obus[temp_w*3 +:temp_w];
assign v226ibus[data_w*3 +:data_w] = c611obus[data_w*0 +:data_w];
assign c611ibus[temp_w*1 +:temp_w] = v376obus[temp_w*1 +:temp_w];
assign v376ibus[data_w*1 +:data_w] = c611obus[data_w*1 +:data_w];
assign c611ibus[temp_w*2 +:temp_w] = v913obus[temp_w*3 +:temp_w];
assign v913ibus[data_w*3 +:data_w] = c611obus[data_w*2 +:data_w];
assign c611ibus[temp_w*3 +:temp_w] = v1013obus[temp_w*1 +:temp_w];
assign v1013ibus[data_w*1 +:data_w] = c611obus[data_w*3 +:data_w];
assign c611ibus[temp_w*4 +:temp_w] = v1763obus[temp_w*1 +:temp_w];
assign v1763ibus[data_w*1 +:data_w] = c611obus[data_w*4 +:data_w];
assign c611ibus[temp_w*5 +:temp_w] = v1859obus[temp_w*0 +:temp_w];
assign v1859ibus[data_w*0 +:data_w] = c611obus[data_w*5 +:data_w];
assign c612ibus[temp_w*0 +:temp_w] = v227obus[temp_w*3 +:temp_w];
assign v227ibus[data_w*3 +:data_w] = c612obus[data_w*0 +:data_w];
assign c612ibus[temp_w*1 +:temp_w] = v377obus[temp_w*1 +:temp_w];
assign v377ibus[data_w*1 +:data_w] = c612obus[data_w*1 +:data_w];
assign c612ibus[temp_w*2 +:temp_w] = v914obus[temp_w*3 +:temp_w];
assign v914ibus[data_w*3 +:data_w] = c612obus[data_w*2 +:data_w];
assign c612ibus[temp_w*3 +:temp_w] = v1014obus[temp_w*1 +:temp_w];
assign v1014ibus[data_w*1 +:data_w] = c612obus[data_w*3 +:data_w];
assign c612ibus[temp_w*4 +:temp_w] = v1764obus[temp_w*1 +:temp_w];
assign v1764ibus[data_w*1 +:data_w] = c612obus[data_w*4 +:data_w];
assign c612ibus[temp_w*5 +:temp_w] = v1860obus[temp_w*0 +:temp_w];
assign v1860ibus[data_w*0 +:data_w] = c612obus[data_w*5 +:data_w];
assign c613ibus[temp_w*0 +:temp_w] = v228obus[temp_w*3 +:temp_w];
assign v228ibus[data_w*3 +:data_w] = c613obus[data_w*0 +:data_w];
assign c613ibus[temp_w*1 +:temp_w] = v378obus[temp_w*1 +:temp_w];
assign v378ibus[data_w*1 +:data_w] = c613obus[data_w*1 +:data_w];
assign c613ibus[temp_w*2 +:temp_w] = v915obus[temp_w*3 +:temp_w];
assign v915ibus[data_w*3 +:data_w] = c613obus[data_w*2 +:data_w];
assign c613ibus[temp_w*3 +:temp_w] = v1015obus[temp_w*1 +:temp_w];
assign v1015ibus[data_w*1 +:data_w] = c613obus[data_w*3 +:data_w];
assign c613ibus[temp_w*4 +:temp_w] = v1765obus[temp_w*1 +:temp_w];
assign v1765ibus[data_w*1 +:data_w] = c613obus[data_w*4 +:data_w];
assign c613ibus[temp_w*5 +:temp_w] = v1861obus[temp_w*0 +:temp_w];
assign v1861ibus[data_w*0 +:data_w] = c613obus[data_w*5 +:data_w];
assign c614ibus[temp_w*0 +:temp_w] = v229obus[temp_w*3 +:temp_w];
assign v229ibus[data_w*3 +:data_w] = c614obus[data_w*0 +:data_w];
assign c614ibus[temp_w*1 +:temp_w] = v379obus[temp_w*1 +:temp_w];
assign v379ibus[data_w*1 +:data_w] = c614obus[data_w*1 +:data_w];
assign c614ibus[temp_w*2 +:temp_w] = v916obus[temp_w*3 +:temp_w];
assign v916ibus[data_w*3 +:data_w] = c614obus[data_w*2 +:data_w];
assign c614ibus[temp_w*3 +:temp_w] = v1016obus[temp_w*1 +:temp_w];
assign v1016ibus[data_w*1 +:data_w] = c614obus[data_w*3 +:data_w];
assign c614ibus[temp_w*4 +:temp_w] = v1766obus[temp_w*1 +:temp_w];
assign v1766ibus[data_w*1 +:data_w] = c614obus[data_w*4 +:data_w];
assign c614ibus[temp_w*5 +:temp_w] = v1862obus[temp_w*0 +:temp_w];
assign v1862ibus[data_w*0 +:data_w] = c614obus[data_w*5 +:data_w];
assign c615ibus[temp_w*0 +:temp_w] = v230obus[temp_w*3 +:temp_w];
assign v230ibus[data_w*3 +:data_w] = c615obus[data_w*0 +:data_w];
assign c615ibus[temp_w*1 +:temp_w] = v380obus[temp_w*1 +:temp_w];
assign v380ibus[data_w*1 +:data_w] = c615obus[data_w*1 +:data_w];
assign c615ibus[temp_w*2 +:temp_w] = v917obus[temp_w*3 +:temp_w];
assign v917ibus[data_w*3 +:data_w] = c615obus[data_w*2 +:data_w];
assign c615ibus[temp_w*3 +:temp_w] = v1017obus[temp_w*1 +:temp_w];
assign v1017ibus[data_w*1 +:data_w] = c615obus[data_w*3 +:data_w];
assign c615ibus[temp_w*4 +:temp_w] = v1767obus[temp_w*1 +:temp_w];
assign v1767ibus[data_w*1 +:data_w] = c615obus[data_w*4 +:data_w];
assign c615ibus[temp_w*5 +:temp_w] = v1863obus[temp_w*0 +:temp_w];
assign v1863ibus[data_w*0 +:data_w] = c615obus[data_w*5 +:data_w];
assign c616ibus[temp_w*0 +:temp_w] = v231obus[temp_w*3 +:temp_w];
assign v231ibus[data_w*3 +:data_w] = c616obus[data_w*0 +:data_w];
assign c616ibus[temp_w*1 +:temp_w] = v381obus[temp_w*1 +:temp_w];
assign v381ibus[data_w*1 +:data_w] = c616obus[data_w*1 +:data_w];
assign c616ibus[temp_w*2 +:temp_w] = v918obus[temp_w*3 +:temp_w];
assign v918ibus[data_w*3 +:data_w] = c616obus[data_w*2 +:data_w];
assign c616ibus[temp_w*3 +:temp_w] = v1018obus[temp_w*1 +:temp_w];
assign v1018ibus[data_w*1 +:data_w] = c616obus[data_w*3 +:data_w];
assign c616ibus[temp_w*4 +:temp_w] = v1768obus[temp_w*1 +:temp_w];
assign v1768ibus[data_w*1 +:data_w] = c616obus[data_w*4 +:data_w];
assign c616ibus[temp_w*5 +:temp_w] = v1864obus[temp_w*0 +:temp_w];
assign v1864ibus[data_w*0 +:data_w] = c616obus[data_w*5 +:data_w];
assign c617ibus[temp_w*0 +:temp_w] = v232obus[temp_w*3 +:temp_w];
assign v232ibus[data_w*3 +:data_w] = c617obus[data_w*0 +:data_w];
assign c617ibus[temp_w*1 +:temp_w] = v382obus[temp_w*1 +:temp_w];
assign v382ibus[data_w*1 +:data_w] = c617obus[data_w*1 +:data_w];
assign c617ibus[temp_w*2 +:temp_w] = v919obus[temp_w*3 +:temp_w];
assign v919ibus[data_w*3 +:data_w] = c617obus[data_w*2 +:data_w];
assign c617ibus[temp_w*3 +:temp_w] = v1019obus[temp_w*1 +:temp_w];
assign v1019ibus[data_w*1 +:data_w] = c617obus[data_w*3 +:data_w];
assign c617ibus[temp_w*4 +:temp_w] = v1769obus[temp_w*1 +:temp_w];
assign v1769ibus[data_w*1 +:data_w] = c617obus[data_w*4 +:data_w];
assign c617ibus[temp_w*5 +:temp_w] = v1865obus[temp_w*0 +:temp_w];
assign v1865ibus[data_w*0 +:data_w] = c617obus[data_w*5 +:data_w];
assign c618ibus[temp_w*0 +:temp_w] = v233obus[temp_w*3 +:temp_w];
assign v233ibus[data_w*3 +:data_w] = c618obus[data_w*0 +:data_w];
assign c618ibus[temp_w*1 +:temp_w] = v383obus[temp_w*1 +:temp_w];
assign v383ibus[data_w*1 +:data_w] = c618obus[data_w*1 +:data_w];
assign c618ibus[temp_w*2 +:temp_w] = v920obus[temp_w*3 +:temp_w];
assign v920ibus[data_w*3 +:data_w] = c618obus[data_w*2 +:data_w];
assign c618ibus[temp_w*3 +:temp_w] = v1020obus[temp_w*1 +:temp_w];
assign v1020ibus[data_w*1 +:data_w] = c618obus[data_w*3 +:data_w];
assign c618ibus[temp_w*4 +:temp_w] = v1770obus[temp_w*1 +:temp_w];
assign v1770ibus[data_w*1 +:data_w] = c618obus[data_w*4 +:data_w];
assign c618ibus[temp_w*5 +:temp_w] = v1866obus[temp_w*0 +:temp_w];
assign v1866ibus[data_w*0 +:data_w] = c618obus[data_w*5 +:data_w];
assign c619ibus[temp_w*0 +:temp_w] = v234obus[temp_w*3 +:temp_w];
assign v234ibus[data_w*3 +:data_w] = c619obus[data_w*0 +:data_w];
assign c619ibus[temp_w*1 +:temp_w] = v288obus[temp_w*1 +:temp_w];
assign v288ibus[data_w*1 +:data_w] = c619obus[data_w*1 +:data_w];
assign c619ibus[temp_w*2 +:temp_w] = v921obus[temp_w*3 +:temp_w];
assign v921ibus[data_w*3 +:data_w] = c619obus[data_w*2 +:data_w];
assign c619ibus[temp_w*3 +:temp_w] = v1021obus[temp_w*1 +:temp_w];
assign v1021ibus[data_w*1 +:data_w] = c619obus[data_w*3 +:data_w];
assign c619ibus[temp_w*4 +:temp_w] = v1771obus[temp_w*1 +:temp_w];
assign v1771ibus[data_w*1 +:data_w] = c619obus[data_w*4 +:data_w];
assign c619ibus[temp_w*5 +:temp_w] = v1867obus[temp_w*0 +:temp_w];
assign v1867ibus[data_w*0 +:data_w] = c619obus[data_w*5 +:data_w];
assign c620ibus[temp_w*0 +:temp_w] = v235obus[temp_w*3 +:temp_w];
assign v235ibus[data_w*3 +:data_w] = c620obus[data_w*0 +:data_w];
assign c620ibus[temp_w*1 +:temp_w] = v289obus[temp_w*1 +:temp_w];
assign v289ibus[data_w*1 +:data_w] = c620obus[data_w*1 +:data_w];
assign c620ibus[temp_w*2 +:temp_w] = v922obus[temp_w*3 +:temp_w];
assign v922ibus[data_w*3 +:data_w] = c620obus[data_w*2 +:data_w];
assign c620ibus[temp_w*3 +:temp_w] = v1022obus[temp_w*1 +:temp_w];
assign v1022ibus[data_w*1 +:data_w] = c620obus[data_w*3 +:data_w];
assign c620ibus[temp_w*4 +:temp_w] = v1772obus[temp_w*1 +:temp_w];
assign v1772ibus[data_w*1 +:data_w] = c620obus[data_w*4 +:data_w];
assign c620ibus[temp_w*5 +:temp_w] = v1868obus[temp_w*0 +:temp_w];
assign v1868ibus[data_w*0 +:data_w] = c620obus[data_w*5 +:data_w];
assign c621ibus[temp_w*0 +:temp_w] = v236obus[temp_w*3 +:temp_w];
assign v236ibus[data_w*3 +:data_w] = c621obus[data_w*0 +:data_w];
assign c621ibus[temp_w*1 +:temp_w] = v290obus[temp_w*1 +:temp_w];
assign v290ibus[data_w*1 +:data_w] = c621obus[data_w*1 +:data_w];
assign c621ibus[temp_w*2 +:temp_w] = v923obus[temp_w*3 +:temp_w];
assign v923ibus[data_w*3 +:data_w] = c621obus[data_w*2 +:data_w];
assign c621ibus[temp_w*3 +:temp_w] = v1023obus[temp_w*1 +:temp_w];
assign v1023ibus[data_w*1 +:data_w] = c621obus[data_w*3 +:data_w];
assign c621ibus[temp_w*4 +:temp_w] = v1773obus[temp_w*1 +:temp_w];
assign v1773ibus[data_w*1 +:data_w] = c621obus[data_w*4 +:data_w];
assign c621ibus[temp_w*5 +:temp_w] = v1869obus[temp_w*0 +:temp_w];
assign v1869ibus[data_w*0 +:data_w] = c621obus[data_w*5 +:data_w];
assign c622ibus[temp_w*0 +:temp_w] = v237obus[temp_w*3 +:temp_w];
assign v237ibus[data_w*3 +:data_w] = c622obus[data_w*0 +:data_w];
assign c622ibus[temp_w*1 +:temp_w] = v291obus[temp_w*1 +:temp_w];
assign v291ibus[data_w*1 +:data_w] = c622obus[data_w*1 +:data_w];
assign c622ibus[temp_w*2 +:temp_w] = v924obus[temp_w*3 +:temp_w];
assign v924ibus[data_w*3 +:data_w] = c622obus[data_w*2 +:data_w];
assign c622ibus[temp_w*3 +:temp_w] = v1024obus[temp_w*1 +:temp_w];
assign v1024ibus[data_w*1 +:data_w] = c622obus[data_w*3 +:data_w];
assign c622ibus[temp_w*4 +:temp_w] = v1774obus[temp_w*1 +:temp_w];
assign v1774ibus[data_w*1 +:data_w] = c622obus[data_w*4 +:data_w];
assign c622ibus[temp_w*5 +:temp_w] = v1870obus[temp_w*0 +:temp_w];
assign v1870ibus[data_w*0 +:data_w] = c622obus[data_w*5 +:data_w];
assign c623ibus[temp_w*0 +:temp_w] = v238obus[temp_w*3 +:temp_w];
assign v238ibus[data_w*3 +:data_w] = c623obus[data_w*0 +:data_w];
assign c623ibus[temp_w*1 +:temp_w] = v292obus[temp_w*1 +:temp_w];
assign v292ibus[data_w*1 +:data_w] = c623obus[data_w*1 +:data_w];
assign c623ibus[temp_w*2 +:temp_w] = v925obus[temp_w*3 +:temp_w];
assign v925ibus[data_w*3 +:data_w] = c623obus[data_w*2 +:data_w];
assign c623ibus[temp_w*3 +:temp_w] = v1025obus[temp_w*1 +:temp_w];
assign v1025ibus[data_w*1 +:data_w] = c623obus[data_w*3 +:data_w];
assign c623ibus[temp_w*4 +:temp_w] = v1775obus[temp_w*1 +:temp_w];
assign v1775ibus[data_w*1 +:data_w] = c623obus[data_w*4 +:data_w];
assign c623ibus[temp_w*5 +:temp_w] = v1871obus[temp_w*0 +:temp_w];
assign v1871ibus[data_w*0 +:data_w] = c623obus[data_w*5 +:data_w];
assign c624ibus[temp_w*0 +:temp_w] = v239obus[temp_w*3 +:temp_w];
assign v239ibus[data_w*3 +:data_w] = c624obus[data_w*0 +:data_w];
assign c624ibus[temp_w*1 +:temp_w] = v293obus[temp_w*1 +:temp_w];
assign v293ibus[data_w*1 +:data_w] = c624obus[data_w*1 +:data_w];
assign c624ibus[temp_w*2 +:temp_w] = v926obus[temp_w*3 +:temp_w];
assign v926ibus[data_w*3 +:data_w] = c624obus[data_w*2 +:data_w];
assign c624ibus[temp_w*3 +:temp_w] = v1026obus[temp_w*1 +:temp_w];
assign v1026ibus[data_w*1 +:data_w] = c624obus[data_w*3 +:data_w];
assign c624ibus[temp_w*4 +:temp_w] = v1776obus[temp_w*1 +:temp_w];
assign v1776ibus[data_w*1 +:data_w] = c624obus[data_w*4 +:data_w];
assign c624ibus[temp_w*5 +:temp_w] = v1872obus[temp_w*0 +:temp_w];
assign v1872ibus[data_w*0 +:data_w] = c624obus[data_w*5 +:data_w];
assign c625ibus[temp_w*0 +:temp_w] = v240obus[temp_w*3 +:temp_w];
assign v240ibus[data_w*3 +:data_w] = c625obus[data_w*0 +:data_w];
assign c625ibus[temp_w*1 +:temp_w] = v294obus[temp_w*1 +:temp_w];
assign v294ibus[data_w*1 +:data_w] = c625obus[data_w*1 +:data_w];
assign c625ibus[temp_w*2 +:temp_w] = v927obus[temp_w*3 +:temp_w];
assign v927ibus[data_w*3 +:data_w] = c625obus[data_w*2 +:data_w];
assign c625ibus[temp_w*3 +:temp_w] = v1027obus[temp_w*1 +:temp_w];
assign v1027ibus[data_w*1 +:data_w] = c625obus[data_w*3 +:data_w];
assign c625ibus[temp_w*4 +:temp_w] = v1777obus[temp_w*1 +:temp_w];
assign v1777ibus[data_w*1 +:data_w] = c625obus[data_w*4 +:data_w];
assign c625ibus[temp_w*5 +:temp_w] = v1873obus[temp_w*0 +:temp_w];
assign v1873ibus[data_w*0 +:data_w] = c625obus[data_w*5 +:data_w];
assign c626ibus[temp_w*0 +:temp_w] = v241obus[temp_w*3 +:temp_w];
assign v241ibus[data_w*3 +:data_w] = c626obus[data_w*0 +:data_w];
assign c626ibus[temp_w*1 +:temp_w] = v295obus[temp_w*1 +:temp_w];
assign v295ibus[data_w*1 +:data_w] = c626obus[data_w*1 +:data_w];
assign c626ibus[temp_w*2 +:temp_w] = v928obus[temp_w*3 +:temp_w];
assign v928ibus[data_w*3 +:data_w] = c626obus[data_w*2 +:data_w];
assign c626ibus[temp_w*3 +:temp_w] = v1028obus[temp_w*1 +:temp_w];
assign v1028ibus[data_w*1 +:data_w] = c626obus[data_w*3 +:data_w];
assign c626ibus[temp_w*4 +:temp_w] = v1778obus[temp_w*1 +:temp_w];
assign v1778ibus[data_w*1 +:data_w] = c626obus[data_w*4 +:data_w];
assign c626ibus[temp_w*5 +:temp_w] = v1874obus[temp_w*0 +:temp_w];
assign v1874ibus[data_w*0 +:data_w] = c626obus[data_w*5 +:data_w];
assign c627ibus[temp_w*0 +:temp_w] = v242obus[temp_w*3 +:temp_w];
assign v242ibus[data_w*3 +:data_w] = c627obus[data_w*0 +:data_w];
assign c627ibus[temp_w*1 +:temp_w] = v296obus[temp_w*1 +:temp_w];
assign v296ibus[data_w*1 +:data_w] = c627obus[data_w*1 +:data_w];
assign c627ibus[temp_w*2 +:temp_w] = v929obus[temp_w*3 +:temp_w];
assign v929ibus[data_w*3 +:data_w] = c627obus[data_w*2 +:data_w];
assign c627ibus[temp_w*3 +:temp_w] = v1029obus[temp_w*1 +:temp_w];
assign v1029ibus[data_w*1 +:data_w] = c627obus[data_w*3 +:data_w];
assign c627ibus[temp_w*4 +:temp_w] = v1779obus[temp_w*1 +:temp_w];
assign v1779ibus[data_w*1 +:data_w] = c627obus[data_w*4 +:data_w];
assign c627ibus[temp_w*5 +:temp_w] = v1875obus[temp_w*0 +:temp_w];
assign v1875ibus[data_w*0 +:data_w] = c627obus[data_w*5 +:data_w];
assign c628ibus[temp_w*0 +:temp_w] = v243obus[temp_w*3 +:temp_w];
assign v243ibus[data_w*3 +:data_w] = c628obus[data_w*0 +:data_w];
assign c628ibus[temp_w*1 +:temp_w] = v297obus[temp_w*1 +:temp_w];
assign v297ibus[data_w*1 +:data_w] = c628obus[data_w*1 +:data_w];
assign c628ibus[temp_w*2 +:temp_w] = v930obus[temp_w*3 +:temp_w];
assign v930ibus[data_w*3 +:data_w] = c628obus[data_w*2 +:data_w];
assign c628ibus[temp_w*3 +:temp_w] = v1030obus[temp_w*1 +:temp_w];
assign v1030ibus[data_w*1 +:data_w] = c628obus[data_w*3 +:data_w];
assign c628ibus[temp_w*4 +:temp_w] = v1780obus[temp_w*1 +:temp_w];
assign v1780ibus[data_w*1 +:data_w] = c628obus[data_w*4 +:data_w];
assign c628ibus[temp_w*5 +:temp_w] = v1876obus[temp_w*0 +:temp_w];
assign v1876ibus[data_w*0 +:data_w] = c628obus[data_w*5 +:data_w];
assign c629ibus[temp_w*0 +:temp_w] = v244obus[temp_w*3 +:temp_w];
assign v244ibus[data_w*3 +:data_w] = c629obus[data_w*0 +:data_w];
assign c629ibus[temp_w*1 +:temp_w] = v298obus[temp_w*1 +:temp_w];
assign v298ibus[data_w*1 +:data_w] = c629obus[data_w*1 +:data_w];
assign c629ibus[temp_w*2 +:temp_w] = v931obus[temp_w*3 +:temp_w];
assign v931ibus[data_w*3 +:data_w] = c629obus[data_w*2 +:data_w];
assign c629ibus[temp_w*3 +:temp_w] = v1031obus[temp_w*1 +:temp_w];
assign v1031ibus[data_w*1 +:data_w] = c629obus[data_w*3 +:data_w];
assign c629ibus[temp_w*4 +:temp_w] = v1781obus[temp_w*1 +:temp_w];
assign v1781ibus[data_w*1 +:data_w] = c629obus[data_w*4 +:data_w];
assign c629ibus[temp_w*5 +:temp_w] = v1877obus[temp_w*0 +:temp_w];
assign v1877ibus[data_w*0 +:data_w] = c629obus[data_w*5 +:data_w];
assign c630ibus[temp_w*0 +:temp_w] = v245obus[temp_w*3 +:temp_w];
assign v245ibus[data_w*3 +:data_w] = c630obus[data_w*0 +:data_w];
assign c630ibus[temp_w*1 +:temp_w] = v299obus[temp_w*1 +:temp_w];
assign v299ibus[data_w*1 +:data_w] = c630obus[data_w*1 +:data_w];
assign c630ibus[temp_w*2 +:temp_w] = v932obus[temp_w*3 +:temp_w];
assign v932ibus[data_w*3 +:data_w] = c630obus[data_w*2 +:data_w];
assign c630ibus[temp_w*3 +:temp_w] = v1032obus[temp_w*1 +:temp_w];
assign v1032ibus[data_w*1 +:data_w] = c630obus[data_w*3 +:data_w];
assign c630ibus[temp_w*4 +:temp_w] = v1782obus[temp_w*1 +:temp_w];
assign v1782ibus[data_w*1 +:data_w] = c630obus[data_w*4 +:data_w];
assign c630ibus[temp_w*5 +:temp_w] = v1878obus[temp_w*0 +:temp_w];
assign v1878ibus[data_w*0 +:data_w] = c630obus[data_w*5 +:data_w];
assign c631ibus[temp_w*0 +:temp_w] = v246obus[temp_w*3 +:temp_w];
assign v246ibus[data_w*3 +:data_w] = c631obus[data_w*0 +:data_w];
assign c631ibus[temp_w*1 +:temp_w] = v300obus[temp_w*1 +:temp_w];
assign v300ibus[data_w*1 +:data_w] = c631obus[data_w*1 +:data_w];
assign c631ibus[temp_w*2 +:temp_w] = v933obus[temp_w*3 +:temp_w];
assign v933ibus[data_w*3 +:data_w] = c631obus[data_w*2 +:data_w];
assign c631ibus[temp_w*3 +:temp_w] = v1033obus[temp_w*1 +:temp_w];
assign v1033ibus[data_w*1 +:data_w] = c631obus[data_w*3 +:data_w];
assign c631ibus[temp_w*4 +:temp_w] = v1783obus[temp_w*1 +:temp_w];
assign v1783ibus[data_w*1 +:data_w] = c631obus[data_w*4 +:data_w];
assign c631ibus[temp_w*5 +:temp_w] = v1879obus[temp_w*0 +:temp_w];
assign v1879ibus[data_w*0 +:data_w] = c631obus[data_w*5 +:data_w];
assign c632ibus[temp_w*0 +:temp_w] = v247obus[temp_w*3 +:temp_w];
assign v247ibus[data_w*3 +:data_w] = c632obus[data_w*0 +:data_w];
assign c632ibus[temp_w*1 +:temp_w] = v301obus[temp_w*1 +:temp_w];
assign v301ibus[data_w*1 +:data_w] = c632obus[data_w*1 +:data_w];
assign c632ibus[temp_w*2 +:temp_w] = v934obus[temp_w*3 +:temp_w];
assign v934ibus[data_w*3 +:data_w] = c632obus[data_w*2 +:data_w];
assign c632ibus[temp_w*3 +:temp_w] = v1034obus[temp_w*1 +:temp_w];
assign v1034ibus[data_w*1 +:data_w] = c632obus[data_w*3 +:data_w];
assign c632ibus[temp_w*4 +:temp_w] = v1784obus[temp_w*1 +:temp_w];
assign v1784ibus[data_w*1 +:data_w] = c632obus[data_w*4 +:data_w];
assign c632ibus[temp_w*5 +:temp_w] = v1880obus[temp_w*0 +:temp_w];
assign v1880ibus[data_w*0 +:data_w] = c632obus[data_w*5 +:data_w];
assign c633ibus[temp_w*0 +:temp_w] = v248obus[temp_w*3 +:temp_w];
assign v248ibus[data_w*3 +:data_w] = c633obus[data_w*0 +:data_w];
assign c633ibus[temp_w*1 +:temp_w] = v302obus[temp_w*1 +:temp_w];
assign v302ibus[data_w*1 +:data_w] = c633obus[data_w*1 +:data_w];
assign c633ibus[temp_w*2 +:temp_w] = v935obus[temp_w*3 +:temp_w];
assign v935ibus[data_w*3 +:data_w] = c633obus[data_w*2 +:data_w];
assign c633ibus[temp_w*3 +:temp_w] = v1035obus[temp_w*1 +:temp_w];
assign v1035ibus[data_w*1 +:data_w] = c633obus[data_w*3 +:data_w];
assign c633ibus[temp_w*4 +:temp_w] = v1785obus[temp_w*1 +:temp_w];
assign v1785ibus[data_w*1 +:data_w] = c633obus[data_w*4 +:data_w];
assign c633ibus[temp_w*5 +:temp_w] = v1881obus[temp_w*0 +:temp_w];
assign v1881ibus[data_w*0 +:data_w] = c633obus[data_w*5 +:data_w];
assign c634ibus[temp_w*0 +:temp_w] = v249obus[temp_w*3 +:temp_w];
assign v249ibus[data_w*3 +:data_w] = c634obus[data_w*0 +:data_w];
assign c634ibus[temp_w*1 +:temp_w] = v303obus[temp_w*1 +:temp_w];
assign v303ibus[data_w*1 +:data_w] = c634obus[data_w*1 +:data_w];
assign c634ibus[temp_w*2 +:temp_w] = v936obus[temp_w*3 +:temp_w];
assign v936ibus[data_w*3 +:data_w] = c634obus[data_w*2 +:data_w];
assign c634ibus[temp_w*3 +:temp_w] = v1036obus[temp_w*1 +:temp_w];
assign v1036ibus[data_w*1 +:data_w] = c634obus[data_w*3 +:data_w];
assign c634ibus[temp_w*4 +:temp_w] = v1786obus[temp_w*1 +:temp_w];
assign v1786ibus[data_w*1 +:data_w] = c634obus[data_w*4 +:data_w];
assign c634ibus[temp_w*5 +:temp_w] = v1882obus[temp_w*0 +:temp_w];
assign v1882ibus[data_w*0 +:data_w] = c634obus[data_w*5 +:data_w];
assign c635ibus[temp_w*0 +:temp_w] = v250obus[temp_w*3 +:temp_w];
assign v250ibus[data_w*3 +:data_w] = c635obus[data_w*0 +:data_w];
assign c635ibus[temp_w*1 +:temp_w] = v304obus[temp_w*1 +:temp_w];
assign v304ibus[data_w*1 +:data_w] = c635obus[data_w*1 +:data_w];
assign c635ibus[temp_w*2 +:temp_w] = v937obus[temp_w*3 +:temp_w];
assign v937ibus[data_w*3 +:data_w] = c635obus[data_w*2 +:data_w];
assign c635ibus[temp_w*3 +:temp_w] = v1037obus[temp_w*1 +:temp_w];
assign v1037ibus[data_w*1 +:data_w] = c635obus[data_w*3 +:data_w];
assign c635ibus[temp_w*4 +:temp_w] = v1787obus[temp_w*1 +:temp_w];
assign v1787ibus[data_w*1 +:data_w] = c635obus[data_w*4 +:data_w];
assign c635ibus[temp_w*5 +:temp_w] = v1883obus[temp_w*0 +:temp_w];
assign v1883ibus[data_w*0 +:data_w] = c635obus[data_w*5 +:data_w];
assign c636ibus[temp_w*0 +:temp_w] = v251obus[temp_w*3 +:temp_w];
assign v251ibus[data_w*3 +:data_w] = c636obus[data_w*0 +:data_w];
assign c636ibus[temp_w*1 +:temp_w] = v305obus[temp_w*1 +:temp_w];
assign v305ibus[data_w*1 +:data_w] = c636obus[data_w*1 +:data_w];
assign c636ibus[temp_w*2 +:temp_w] = v938obus[temp_w*3 +:temp_w];
assign v938ibus[data_w*3 +:data_w] = c636obus[data_w*2 +:data_w];
assign c636ibus[temp_w*3 +:temp_w] = v1038obus[temp_w*1 +:temp_w];
assign v1038ibus[data_w*1 +:data_w] = c636obus[data_w*3 +:data_w];
assign c636ibus[temp_w*4 +:temp_w] = v1788obus[temp_w*1 +:temp_w];
assign v1788ibus[data_w*1 +:data_w] = c636obus[data_w*4 +:data_w];
assign c636ibus[temp_w*5 +:temp_w] = v1884obus[temp_w*0 +:temp_w];
assign v1884ibus[data_w*0 +:data_w] = c636obus[data_w*5 +:data_w];
assign c637ibus[temp_w*0 +:temp_w] = v252obus[temp_w*3 +:temp_w];
assign v252ibus[data_w*3 +:data_w] = c637obus[data_w*0 +:data_w];
assign c637ibus[temp_w*1 +:temp_w] = v306obus[temp_w*1 +:temp_w];
assign v306ibus[data_w*1 +:data_w] = c637obus[data_w*1 +:data_w];
assign c637ibus[temp_w*2 +:temp_w] = v939obus[temp_w*3 +:temp_w];
assign v939ibus[data_w*3 +:data_w] = c637obus[data_w*2 +:data_w];
assign c637ibus[temp_w*3 +:temp_w] = v1039obus[temp_w*1 +:temp_w];
assign v1039ibus[data_w*1 +:data_w] = c637obus[data_w*3 +:data_w];
assign c637ibus[temp_w*4 +:temp_w] = v1789obus[temp_w*1 +:temp_w];
assign v1789ibus[data_w*1 +:data_w] = c637obus[data_w*4 +:data_w];
assign c637ibus[temp_w*5 +:temp_w] = v1885obus[temp_w*0 +:temp_w];
assign v1885ibus[data_w*0 +:data_w] = c637obus[data_w*5 +:data_w];
assign c638ibus[temp_w*0 +:temp_w] = v253obus[temp_w*3 +:temp_w];
assign v253ibus[data_w*3 +:data_w] = c638obus[data_w*0 +:data_w];
assign c638ibus[temp_w*1 +:temp_w] = v307obus[temp_w*1 +:temp_w];
assign v307ibus[data_w*1 +:data_w] = c638obus[data_w*1 +:data_w];
assign c638ibus[temp_w*2 +:temp_w] = v940obus[temp_w*3 +:temp_w];
assign v940ibus[data_w*3 +:data_w] = c638obus[data_w*2 +:data_w];
assign c638ibus[temp_w*3 +:temp_w] = v1040obus[temp_w*1 +:temp_w];
assign v1040ibus[data_w*1 +:data_w] = c638obus[data_w*3 +:data_w];
assign c638ibus[temp_w*4 +:temp_w] = v1790obus[temp_w*1 +:temp_w];
assign v1790ibus[data_w*1 +:data_w] = c638obus[data_w*4 +:data_w];
assign c638ibus[temp_w*5 +:temp_w] = v1886obus[temp_w*0 +:temp_w];
assign v1886ibus[data_w*0 +:data_w] = c638obus[data_w*5 +:data_w];
assign c639ibus[temp_w*0 +:temp_w] = v254obus[temp_w*3 +:temp_w];
assign v254ibus[data_w*3 +:data_w] = c639obus[data_w*0 +:data_w];
assign c639ibus[temp_w*1 +:temp_w] = v308obus[temp_w*1 +:temp_w];
assign v308ibus[data_w*1 +:data_w] = c639obus[data_w*1 +:data_w];
assign c639ibus[temp_w*2 +:temp_w] = v941obus[temp_w*3 +:temp_w];
assign v941ibus[data_w*3 +:data_w] = c639obus[data_w*2 +:data_w];
assign c639ibus[temp_w*3 +:temp_w] = v1041obus[temp_w*1 +:temp_w];
assign v1041ibus[data_w*1 +:data_w] = c639obus[data_w*3 +:data_w];
assign c639ibus[temp_w*4 +:temp_w] = v1791obus[temp_w*1 +:temp_w];
assign v1791ibus[data_w*1 +:data_w] = c639obus[data_w*4 +:data_w];
assign c639ibus[temp_w*5 +:temp_w] = v1887obus[temp_w*0 +:temp_w];
assign v1887ibus[data_w*0 +:data_w] = c639obus[data_w*5 +:data_w];
assign c640ibus[temp_w*0 +:temp_w] = v255obus[temp_w*3 +:temp_w];
assign v255ibus[data_w*3 +:data_w] = c640obus[data_w*0 +:data_w];
assign c640ibus[temp_w*1 +:temp_w] = v309obus[temp_w*1 +:temp_w];
assign v309ibus[data_w*1 +:data_w] = c640obus[data_w*1 +:data_w];
assign c640ibus[temp_w*2 +:temp_w] = v942obus[temp_w*3 +:temp_w];
assign v942ibus[data_w*3 +:data_w] = c640obus[data_w*2 +:data_w];
assign c640ibus[temp_w*3 +:temp_w] = v1042obus[temp_w*1 +:temp_w];
assign v1042ibus[data_w*1 +:data_w] = c640obus[data_w*3 +:data_w];
assign c640ibus[temp_w*4 +:temp_w] = v1792obus[temp_w*1 +:temp_w];
assign v1792ibus[data_w*1 +:data_w] = c640obus[data_w*4 +:data_w];
assign c640ibus[temp_w*5 +:temp_w] = v1888obus[temp_w*0 +:temp_w];
assign v1888ibus[data_w*0 +:data_w] = c640obus[data_w*5 +:data_w];
assign c641ibus[temp_w*0 +:temp_w] = v256obus[temp_w*3 +:temp_w];
assign v256ibus[data_w*3 +:data_w] = c641obus[data_w*0 +:data_w];
assign c641ibus[temp_w*1 +:temp_w] = v310obus[temp_w*1 +:temp_w];
assign v310ibus[data_w*1 +:data_w] = c641obus[data_w*1 +:data_w];
assign c641ibus[temp_w*2 +:temp_w] = v943obus[temp_w*3 +:temp_w];
assign v943ibus[data_w*3 +:data_w] = c641obus[data_w*2 +:data_w];
assign c641ibus[temp_w*3 +:temp_w] = v1043obus[temp_w*1 +:temp_w];
assign v1043ibus[data_w*1 +:data_w] = c641obus[data_w*3 +:data_w];
assign c641ibus[temp_w*4 +:temp_w] = v1793obus[temp_w*1 +:temp_w];
assign v1793ibus[data_w*1 +:data_w] = c641obus[data_w*4 +:data_w];
assign c641ibus[temp_w*5 +:temp_w] = v1889obus[temp_w*0 +:temp_w];
assign v1889ibus[data_w*0 +:data_w] = c641obus[data_w*5 +:data_w];
assign c642ibus[temp_w*0 +:temp_w] = v257obus[temp_w*3 +:temp_w];
assign v257ibus[data_w*3 +:data_w] = c642obus[data_w*0 +:data_w];
assign c642ibus[temp_w*1 +:temp_w] = v311obus[temp_w*1 +:temp_w];
assign v311ibus[data_w*1 +:data_w] = c642obus[data_w*1 +:data_w];
assign c642ibus[temp_w*2 +:temp_w] = v944obus[temp_w*3 +:temp_w];
assign v944ibus[data_w*3 +:data_w] = c642obus[data_w*2 +:data_w];
assign c642ibus[temp_w*3 +:temp_w] = v1044obus[temp_w*1 +:temp_w];
assign v1044ibus[data_w*1 +:data_w] = c642obus[data_w*3 +:data_w];
assign c642ibus[temp_w*4 +:temp_w] = v1794obus[temp_w*1 +:temp_w];
assign v1794ibus[data_w*1 +:data_w] = c642obus[data_w*4 +:data_w];
assign c642ibus[temp_w*5 +:temp_w] = v1890obus[temp_w*0 +:temp_w];
assign v1890ibus[data_w*0 +:data_w] = c642obus[data_w*5 +:data_w];
assign c643ibus[temp_w*0 +:temp_w] = v258obus[temp_w*3 +:temp_w];
assign v258ibus[data_w*3 +:data_w] = c643obus[data_w*0 +:data_w];
assign c643ibus[temp_w*1 +:temp_w] = v312obus[temp_w*1 +:temp_w];
assign v312ibus[data_w*1 +:data_w] = c643obus[data_w*1 +:data_w];
assign c643ibus[temp_w*2 +:temp_w] = v945obus[temp_w*3 +:temp_w];
assign v945ibus[data_w*3 +:data_w] = c643obus[data_w*2 +:data_w];
assign c643ibus[temp_w*3 +:temp_w] = v1045obus[temp_w*1 +:temp_w];
assign v1045ibus[data_w*1 +:data_w] = c643obus[data_w*3 +:data_w];
assign c643ibus[temp_w*4 +:temp_w] = v1795obus[temp_w*1 +:temp_w];
assign v1795ibus[data_w*1 +:data_w] = c643obus[data_w*4 +:data_w];
assign c643ibus[temp_w*5 +:temp_w] = v1891obus[temp_w*0 +:temp_w];
assign v1891ibus[data_w*0 +:data_w] = c643obus[data_w*5 +:data_w];
assign c644ibus[temp_w*0 +:temp_w] = v259obus[temp_w*3 +:temp_w];
assign v259ibus[data_w*3 +:data_w] = c644obus[data_w*0 +:data_w];
assign c644ibus[temp_w*1 +:temp_w] = v313obus[temp_w*1 +:temp_w];
assign v313ibus[data_w*1 +:data_w] = c644obus[data_w*1 +:data_w];
assign c644ibus[temp_w*2 +:temp_w] = v946obus[temp_w*3 +:temp_w];
assign v946ibus[data_w*3 +:data_w] = c644obus[data_w*2 +:data_w];
assign c644ibus[temp_w*3 +:temp_w] = v1046obus[temp_w*1 +:temp_w];
assign v1046ibus[data_w*1 +:data_w] = c644obus[data_w*3 +:data_w];
assign c644ibus[temp_w*4 +:temp_w] = v1796obus[temp_w*1 +:temp_w];
assign v1796ibus[data_w*1 +:data_w] = c644obus[data_w*4 +:data_w];
assign c644ibus[temp_w*5 +:temp_w] = v1892obus[temp_w*0 +:temp_w];
assign v1892ibus[data_w*0 +:data_w] = c644obus[data_w*5 +:data_w];
assign c645ibus[temp_w*0 +:temp_w] = v260obus[temp_w*3 +:temp_w];
assign v260ibus[data_w*3 +:data_w] = c645obus[data_w*0 +:data_w];
assign c645ibus[temp_w*1 +:temp_w] = v314obus[temp_w*1 +:temp_w];
assign v314ibus[data_w*1 +:data_w] = c645obus[data_w*1 +:data_w];
assign c645ibus[temp_w*2 +:temp_w] = v947obus[temp_w*3 +:temp_w];
assign v947ibus[data_w*3 +:data_w] = c645obus[data_w*2 +:data_w];
assign c645ibus[temp_w*3 +:temp_w] = v1047obus[temp_w*1 +:temp_w];
assign v1047ibus[data_w*1 +:data_w] = c645obus[data_w*3 +:data_w];
assign c645ibus[temp_w*4 +:temp_w] = v1797obus[temp_w*1 +:temp_w];
assign v1797ibus[data_w*1 +:data_w] = c645obus[data_w*4 +:data_w];
assign c645ibus[temp_w*5 +:temp_w] = v1893obus[temp_w*0 +:temp_w];
assign v1893ibus[data_w*0 +:data_w] = c645obus[data_w*5 +:data_w];
assign c646ibus[temp_w*0 +:temp_w] = v261obus[temp_w*3 +:temp_w];
assign v261ibus[data_w*3 +:data_w] = c646obus[data_w*0 +:data_w];
assign c646ibus[temp_w*1 +:temp_w] = v315obus[temp_w*1 +:temp_w];
assign v315ibus[data_w*1 +:data_w] = c646obus[data_w*1 +:data_w];
assign c646ibus[temp_w*2 +:temp_w] = v948obus[temp_w*3 +:temp_w];
assign v948ibus[data_w*3 +:data_w] = c646obus[data_w*2 +:data_w];
assign c646ibus[temp_w*3 +:temp_w] = v1048obus[temp_w*1 +:temp_w];
assign v1048ibus[data_w*1 +:data_w] = c646obus[data_w*3 +:data_w];
assign c646ibus[temp_w*4 +:temp_w] = v1798obus[temp_w*1 +:temp_w];
assign v1798ibus[data_w*1 +:data_w] = c646obus[data_w*4 +:data_w];
assign c646ibus[temp_w*5 +:temp_w] = v1894obus[temp_w*0 +:temp_w];
assign v1894ibus[data_w*0 +:data_w] = c646obus[data_w*5 +:data_w];
assign c647ibus[temp_w*0 +:temp_w] = v262obus[temp_w*3 +:temp_w];
assign v262ibus[data_w*3 +:data_w] = c647obus[data_w*0 +:data_w];
assign c647ibus[temp_w*1 +:temp_w] = v316obus[temp_w*1 +:temp_w];
assign v316ibus[data_w*1 +:data_w] = c647obus[data_w*1 +:data_w];
assign c647ibus[temp_w*2 +:temp_w] = v949obus[temp_w*3 +:temp_w];
assign v949ibus[data_w*3 +:data_w] = c647obus[data_w*2 +:data_w];
assign c647ibus[temp_w*3 +:temp_w] = v1049obus[temp_w*1 +:temp_w];
assign v1049ibus[data_w*1 +:data_w] = c647obus[data_w*3 +:data_w];
assign c647ibus[temp_w*4 +:temp_w] = v1799obus[temp_w*1 +:temp_w];
assign v1799ibus[data_w*1 +:data_w] = c647obus[data_w*4 +:data_w];
assign c647ibus[temp_w*5 +:temp_w] = v1895obus[temp_w*0 +:temp_w];
assign v1895ibus[data_w*0 +:data_w] = c647obus[data_w*5 +:data_w];
assign c648ibus[temp_w*0 +:temp_w] = v263obus[temp_w*3 +:temp_w];
assign v263ibus[data_w*3 +:data_w] = c648obus[data_w*0 +:data_w];
assign c648ibus[temp_w*1 +:temp_w] = v317obus[temp_w*1 +:temp_w];
assign v317ibus[data_w*1 +:data_w] = c648obus[data_w*1 +:data_w];
assign c648ibus[temp_w*2 +:temp_w] = v950obus[temp_w*3 +:temp_w];
assign v950ibus[data_w*3 +:data_w] = c648obus[data_w*2 +:data_w];
assign c648ibus[temp_w*3 +:temp_w] = v1050obus[temp_w*1 +:temp_w];
assign v1050ibus[data_w*1 +:data_w] = c648obus[data_w*3 +:data_w];
assign c648ibus[temp_w*4 +:temp_w] = v1800obus[temp_w*1 +:temp_w];
assign v1800ibus[data_w*1 +:data_w] = c648obus[data_w*4 +:data_w];
assign c648ibus[temp_w*5 +:temp_w] = v1896obus[temp_w*0 +:temp_w];
assign v1896ibus[data_w*0 +:data_w] = c648obus[data_w*5 +:data_w];
assign c649ibus[temp_w*0 +:temp_w] = v264obus[temp_w*3 +:temp_w];
assign v264ibus[data_w*3 +:data_w] = c649obus[data_w*0 +:data_w];
assign c649ibus[temp_w*1 +:temp_w] = v318obus[temp_w*1 +:temp_w];
assign v318ibus[data_w*1 +:data_w] = c649obus[data_w*1 +:data_w];
assign c649ibus[temp_w*2 +:temp_w] = v951obus[temp_w*3 +:temp_w];
assign v951ibus[data_w*3 +:data_w] = c649obus[data_w*2 +:data_w];
assign c649ibus[temp_w*3 +:temp_w] = v1051obus[temp_w*1 +:temp_w];
assign v1051ibus[data_w*1 +:data_w] = c649obus[data_w*3 +:data_w];
assign c649ibus[temp_w*4 +:temp_w] = v1801obus[temp_w*1 +:temp_w];
assign v1801ibus[data_w*1 +:data_w] = c649obus[data_w*4 +:data_w];
assign c649ibus[temp_w*5 +:temp_w] = v1897obus[temp_w*0 +:temp_w];
assign v1897ibus[data_w*0 +:data_w] = c649obus[data_w*5 +:data_w];
assign c650ibus[temp_w*0 +:temp_w] = v265obus[temp_w*3 +:temp_w];
assign v265ibus[data_w*3 +:data_w] = c650obus[data_w*0 +:data_w];
assign c650ibus[temp_w*1 +:temp_w] = v319obus[temp_w*1 +:temp_w];
assign v319ibus[data_w*1 +:data_w] = c650obus[data_w*1 +:data_w];
assign c650ibus[temp_w*2 +:temp_w] = v952obus[temp_w*3 +:temp_w];
assign v952ibus[data_w*3 +:data_w] = c650obus[data_w*2 +:data_w];
assign c650ibus[temp_w*3 +:temp_w] = v1052obus[temp_w*1 +:temp_w];
assign v1052ibus[data_w*1 +:data_w] = c650obus[data_w*3 +:data_w];
assign c650ibus[temp_w*4 +:temp_w] = v1802obus[temp_w*1 +:temp_w];
assign v1802ibus[data_w*1 +:data_w] = c650obus[data_w*4 +:data_w];
assign c650ibus[temp_w*5 +:temp_w] = v1898obus[temp_w*0 +:temp_w];
assign v1898ibus[data_w*0 +:data_w] = c650obus[data_w*5 +:data_w];
assign c651ibus[temp_w*0 +:temp_w] = v266obus[temp_w*3 +:temp_w];
assign v266ibus[data_w*3 +:data_w] = c651obus[data_w*0 +:data_w];
assign c651ibus[temp_w*1 +:temp_w] = v320obus[temp_w*1 +:temp_w];
assign v320ibus[data_w*1 +:data_w] = c651obus[data_w*1 +:data_w];
assign c651ibus[temp_w*2 +:temp_w] = v953obus[temp_w*3 +:temp_w];
assign v953ibus[data_w*3 +:data_w] = c651obus[data_w*2 +:data_w];
assign c651ibus[temp_w*3 +:temp_w] = v1053obus[temp_w*1 +:temp_w];
assign v1053ibus[data_w*1 +:data_w] = c651obus[data_w*3 +:data_w];
assign c651ibus[temp_w*4 +:temp_w] = v1803obus[temp_w*1 +:temp_w];
assign v1803ibus[data_w*1 +:data_w] = c651obus[data_w*4 +:data_w];
assign c651ibus[temp_w*5 +:temp_w] = v1899obus[temp_w*0 +:temp_w];
assign v1899ibus[data_w*0 +:data_w] = c651obus[data_w*5 +:data_w];
assign c652ibus[temp_w*0 +:temp_w] = v267obus[temp_w*3 +:temp_w];
assign v267ibus[data_w*3 +:data_w] = c652obus[data_w*0 +:data_w];
assign c652ibus[temp_w*1 +:temp_w] = v321obus[temp_w*1 +:temp_w];
assign v321ibus[data_w*1 +:data_w] = c652obus[data_w*1 +:data_w];
assign c652ibus[temp_w*2 +:temp_w] = v954obus[temp_w*3 +:temp_w];
assign v954ibus[data_w*3 +:data_w] = c652obus[data_w*2 +:data_w];
assign c652ibus[temp_w*3 +:temp_w] = v1054obus[temp_w*1 +:temp_w];
assign v1054ibus[data_w*1 +:data_w] = c652obus[data_w*3 +:data_w];
assign c652ibus[temp_w*4 +:temp_w] = v1804obus[temp_w*1 +:temp_w];
assign v1804ibus[data_w*1 +:data_w] = c652obus[data_w*4 +:data_w];
assign c652ibus[temp_w*5 +:temp_w] = v1900obus[temp_w*0 +:temp_w];
assign v1900ibus[data_w*0 +:data_w] = c652obus[data_w*5 +:data_w];
assign c653ibus[temp_w*0 +:temp_w] = v268obus[temp_w*3 +:temp_w];
assign v268ibus[data_w*3 +:data_w] = c653obus[data_w*0 +:data_w];
assign c653ibus[temp_w*1 +:temp_w] = v322obus[temp_w*1 +:temp_w];
assign v322ibus[data_w*1 +:data_w] = c653obus[data_w*1 +:data_w];
assign c653ibus[temp_w*2 +:temp_w] = v955obus[temp_w*3 +:temp_w];
assign v955ibus[data_w*3 +:data_w] = c653obus[data_w*2 +:data_w];
assign c653ibus[temp_w*3 +:temp_w] = v1055obus[temp_w*1 +:temp_w];
assign v1055ibus[data_w*1 +:data_w] = c653obus[data_w*3 +:data_w];
assign c653ibus[temp_w*4 +:temp_w] = v1805obus[temp_w*1 +:temp_w];
assign v1805ibus[data_w*1 +:data_w] = c653obus[data_w*4 +:data_w];
assign c653ibus[temp_w*5 +:temp_w] = v1901obus[temp_w*0 +:temp_w];
assign v1901ibus[data_w*0 +:data_w] = c653obus[data_w*5 +:data_w];
assign c654ibus[temp_w*0 +:temp_w] = v269obus[temp_w*3 +:temp_w];
assign v269ibus[data_w*3 +:data_w] = c654obus[data_w*0 +:data_w];
assign c654ibus[temp_w*1 +:temp_w] = v323obus[temp_w*1 +:temp_w];
assign v323ibus[data_w*1 +:data_w] = c654obus[data_w*1 +:data_w];
assign c654ibus[temp_w*2 +:temp_w] = v956obus[temp_w*3 +:temp_w];
assign v956ibus[data_w*3 +:data_w] = c654obus[data_w*2 +:data_w];
assign c654ibus[temp_w*3 +:temp_w] = v960obus[temp_w*1 +:temp_w];
assign v960ibus[data_w*1 +:data_w] = c654obus[data_w*3 +:data_w];
assign c654ibus[temp_w*4 +:temp_w] = v1806obus[temp_w*1 +:temp_w];
assign v1806ibus[data_w*1 +:data_w] = c654obus[data_w*4 +:data_w];
assign c654ibus[temp_w*5 +:temp_w] = v1902obus[temp_w*0 +:temp_w];
assign v1902ibus[data_w*0 +:data_w] = c654obus[data_w*5 +:data_w];
assign c655ibus[temp_w*0 +:temp_w] = v270obus[temp_w*3 +:temp_w];
assign v270ibus[data_w*3 +:data_w] = c655obus[data_w*0 +:data_w];
assign c655ibus[temp_w*1 +:temp_w] = v324obus[temp_w*1 +:temp_w];
assign v324ibus[data_w*1 +:data_w] = c655obus[data_w*1 +:data_w];
assign c655ibus[temp_w*2 +:temp_w] = v957obus[temp_w*3 +:temp_w];
assign v957ibus[data_w*3 +:data_w] = c655obus[data_w*2 +:data_w];
assign c655ibus[temp_w*3 +:temp_w] = v961obus[temp_w*1 +:temp_w];
assign v961ibus[data_w*1 +:data_w] = c655obus[data_w*3 +:data_w];
assign c655ibus[temp_w*4 +:temp_w] = v1807obus[temp_w*1 +:temp_w];
assign v1807ibus[data_w*1 +:data_w] = c655obus[data_w*4 +:data_w];
assign c655ibus[temp_w*5 +:temp_w] = v1903obus[temp_w*0 +:temp_w];
assign v1903ibus[data_w*0 +:data_w] = c655obus[data_w*5 +:data_w];
assign c656ibus[temp_w*0 +:temp_w] = v271obus[temp_w*3 +:temp_w];
assign v271ibus[data_w*3 +:data_w] = c656obus[data_w*0 +:data_w];
assign c656ibus[temp_w*1 +:temp_w] = v325obus[temp_w*1 +:temp_w];
assign v325ibus[data_w*1 +:data_w] = c656obus[data_w*1 +:data_w];
assign c656ibus[temp_w*2 +:temp_w] = v958obus[temp_w*3 +:temp_w];
assign v958ibus[data_w*3 +:data_w] = c656obus[data_w*2 +:data_w];
assign c656ibus[temp_w*3 +:temp_w] = v962obus[temp_w*1 +:temp_w];
assign v962ibus[data_w*1 +:data_w] = c656obus[data_w*3 +:data_w];
assign c656ibus[temp_w*4 +:temp_w] = v1808obus[temp_w*1 +:temp_w];
assign v1808ibus[data_w*1 +:data_w] = c656obus[data_w*4 +:data_w];
assign c656ibus[temp_w*5 +:temp_w] = v1904obus[temp_w*0 +:temp_w];
assign v1904ibus[data_w*0 +:data_w] = c656obus[data_w*5 +:data_w];
assign c657ibus[temp_w*0 +:temp_w] = v272obus[temp_w*3 +:temp_w];
assign v272ibus[data_w*3 +:data_w] = c657obus[data_w*0 +:data_w];
assign c657ibus[temp_w*1 +:temp_w] = v326obus[temp_w*1 +:temp_w];
assign v326ibus[data_w*1 +:data_w] = c657obus[data_w*1 +:data_w];
assign c657ibus[temp_w*2 +:temp_w] = v959obus[temp_w*3 +:temp_w];
assign v959ibus[data_w*3 +:data_w] = c657obus[data_w*2 +:data_w];
assign c657ibus[temp_w*3 +:temp_w] = v963obus[temp_w*1 +:temp_w];
assign v963ibus[data_w*1 +:data_w] = c657obus[data_w*3 +:data_w];
assign c657ibus[temp_w*4 +:temp_w] = v1809obus[temp_w*1 +:temp_w];
assign v1809ibus[data_w*1 +:data_w] = c657obus[data_w*4 +:data_w];
assign c657ibus[temp_w*5 +:temp_w] = v1905obus[temp_w*0 +:temp_w];
assign v1905ibus[data_w*0 +:data_w] = c657obus[data_w*5 +:data_w];
assign c658ibus[temp_w*0 +:temp_w] = v273obus[temp_w*3 +:temp_w];
assign v273ibus[data_w*3 +:data_w] = c658obus[data_w*0 +:data_w];
assign c658ibus[temp_w*1 +:temp_w] = v327obus[temp_w*1 +:temp_w];
assign v327ibus[data_w*1 +:data_w] = c658obus[data_w*1 +:data_w];
assign c658ibus[temp_w*2 +:temp_w] = v864obus[temp_w*3 +:temp_w];
assign v864ibus[data_w*3 +:data_w] = c658obus[data_w*2 +:data_w];
assign c658ibus[temp_w*3 +:temp_w] = v964obus[temp_w*1 +:temp_w];
assign v964ibus[data_w*1 +:data_w] = c658obus[data_w*3 +:data_w];
assign c658ibus[temp_w*4 +:temp_w] = v1810obus[temp_w*1 +:temp_w];
assign v1810ibus[data_w*1 +:data_w] = c658obus[data_w*4 +:data_w];
assign c658ibus[temp_w*5 +:temp_w] = v1906obus[temp_w*0 +:temp_w];
assign v1906ibus[data_w*0 +:data_w] = c658obus[data_w*5 +:data_w];
assign c659ibus[temp_w*0 +:temp_w] = v274obus[temp_w*3 +:temp_w];
assign v274ibus[data_w*3 +:data_w] = c659obus[data_w*0 +:data_w];
assign c659ibus[temp_w*1 +:temp_w] = v328obus[temp_w*1 +:temp_w];
assign v328ibus[data_w*1 +:data_w] = c659obus[data_w*1 +:data_w];
assign c659ibus[temp_w*2 +:temp_w] = v865obus[temp_w*3 +:temp_w];
assign v865ibus[data_w*3 +:data_w] = c659obus[data_w*2 +:data_w];
assign c659ibus[temp_w*3 +:temp_w] = v965obus[temp_w*1 +:temp_w];
assign v965ibus[data_w*1 +:data_w] = c659obus[data_w*3 +:data_w];
assign c659ibus[temp_w*4 +:temp_w] = v1811obus[temp_w*1 +:temp_w];
assign v1811ibus[data_w*1 +:data_w] = c659obus[data_w*4 +:data_w];
assign c659ibus[temp_w*5 +:temp_w] = v1907obus[temp_w*0 +:temp_w];
assign v1907ibus[data_w*0 +:data_w] = c659obus[data_w*5 +:data_w];
assign c660ibus[temp_w*0 +:temp_w] = v275obus[temp_w*3 +:temp_w];
assign v275ibus[data_w*3 +:data_w] = c660obus[data_w*0 +:data_w];
assign c660ibus[temp_w*1 +:temp_w] = v329obus[temp_w*1 +:temp_w];
assign v329ibus[data_w*1 +:data_w] = c660obus[data_w*1 +:data_w];
assign c660ibus[temp_w*2 +:temp_w] = v866obus[temp_w*3 +:temp_w];
assign v866ibus[data_w*3 +:data_w] = c660obus[data_w*2 +:data_w];
assign c660ibus[temp_w*3 +:temp_w] = v966obus[temp_w*1 +:temp_w];
assign v966ibus[data_w*1 +:data_w] = c660obus[data_w*3 +:data_w];
assign c660ibus[temp_w*4 +:temp_w] = v1812obus[temp_w*1 +:temp_w];
assign v1812ibus[data_w*1 +:data_w] = c660obus[data_w*4 +:data_w];
assign c660ibus[temp_w*5 +:temp_w] = v1908obus[temp_w*0 +:temp_w];
assign v1908ibus[data_w*0 +:data_w] = c660obus[data_w*5 +:data_w];
assign c661ibus[temp_w*0 +:temp_w] = v276obus[temp_w*3 +:temp_w];
assign v276ibus[data_w*3 +:data_w] = c661obus[data_w*0 +:data_w];
assign c661ibus[temp_w*1 +:temp_w] = v330obus[temp_w*1 +:temp_w];
assign v330ibus[data_w*1 +:data_w] = c661obus[data_w*1 +:data_w];
assign c661ibus[temp_w*2 +:temp_w] = v867obus[temp_w*3 +:temp_w];
assign v867ibus[data_w*3 +:data_w] = c661obus[data_w*2 +:data_w];
assign c661ibus[temp_w*3 +:temp_w] = v967obus[temp_w*1 +:temp_w];
assign v967ibus[data_w*1 +:data_w] = c661obus[data_w*3 +:data_w];
assign c661ibus[temp_w*4 +:temp_w] = v1813obus[temp_w*1 +:temp_w];
assign v1813ibus[data_w*1 +:data_w] = c661obus[data_w*4 +:data_w];
assign c661ibus[temp_w*5 +:temp_w] = v1909obus[temp_w*0 +:temp_w];
assign v1909ibus[data_w*0 +:data_w] = c661obus[data_w*5 +:data_w];
assign c662ibus[temp_w*0 +:temp_w] = v277obus[temp_w*3 +:temp_w];
assign v277ibus[data_w*3 +:data_w] = c662obus[data_w*0 +:data_w];
assign c662ibus[temp_w*1 +:temp_w] = v331obus[temp_w*1 +:temp_w];
assign v331ibus[data_w*1 +:data_w] = c662obus[data_w*1 +:data_w];
assign c662ibus[temp_w*2 +:temp_w] = v868obus[temp_w*3 +:temp_w];
assign v868ibus[data_w*3 +:data_w] = c662obus[data_w*2 +:data_w];
assign c662ibus[temp_w*3 +:temp_w] = v968obus[temp_w*1 +:temp_w];
assign v968ibus[data_w*1 +:data_w] = c662obus[data_w*3 +:data_w];
assign c662ibus[temp_w*4 +:temp_w] = v1814obus[temp_w*1 +:temp_w];
assign v1814ibus[data_w*1 +:data_w] = c662obus[data_w*4 +:data_w];
assign c662ibus[temp_w*5 +:temp_w] = v1910obus[temp_w*0 +:temp_w];
assign v1910ibus[data_w*0 +:data_w] = c662obus[data_w*5 +:data_w];
assign c663ibus[temp_w*0 +:temp_w] = v278obus[temp_w*3 +:temp_w];
assign v278ibus[data_w*3 +:data_w] = c663obus[data_w*0 +:data_w];
assign c663ibus[temp_w*1 +:temp_w] = v332obus[temp_w*1 +:temp_w];
assign v332ibus[data_w*1 +:data_w] = c663obus[data_w*1 +:data_w];
assign c663ibus[temp_w*2 +:temp_w] = v869obus[temp_w*3 +:temp_w];
assign v869ibus[data_w*3 +:data_w] = c663obus[data_w*2 +:data_w];
assign c663ibus[temp_w*3 +:temp_w] = v969obus[temp_w*1 +:temp_w];
assign v969ibus[data_w*1 +:data_w] = c663obus[data_w*3 +:data_w];
assign c663ibus[temp_w*4 +:temp_w] = v1815obus[temp_w*1 +:temp_w];
assign v1815ibus[data_w*1 +:data_w] = c663obus[data_w*4 +:data_w];
assign c663ibus[temp_w*5 +:temp_w] = v1911obus[temp_w*0 +:temp_w];
assign v1911ibus[data_w*0 +:data_w] = c663obus[data_w*5 +:data_w];
assign c664ibus[temp_w*0 +:temp_w] = v279obus[temp_w*3 +:temp_w];
assign v279ibus[data_w*3 +:data_w] = c664obus[data_w*0 +:data_w];
assign c664ibus[temp_w*1 +:temp_w] = v333obus[temp_w*1 +:temp_w];
assign v333ibus[data_w*1 +:data_w] = c664obus[data_w*1 +:data_w];
assign c664ibus[temp_w*2 +:temp_w] = v870obus[temp_w*3 +:temp_w];
assign v870ibus[data_w*3 +:data_w] = c664obus[data_w*2 +:data_w];
assign c664ibus[temp_w*3 +:temp_w] = v970obus[temp_w*1 +:temp_w];
assign v970ibus[data_w*1 +:data_w] = c664obus[data_w*3 +:data_w];
assign c664ibus[temp_w*4 +:temp_w] = v1816obus[temp_w*1 +:temp_w];
assign v1816ibus[data_w*1 +:data_w] = c664obus[data_w*4 +:data_w];
assign c664ibus[temp_w*5 +:temp_w] = v1912obus[temp_w*0 +:temp_w];
assign v1912ibus[data_w*0 +:data_w] = c664obus[data_w*5 +:data_w];
assign c665ibus[temp_w*0 +:temp_w] = v280obus[temp_w*3 +:temp_w];
assign v280ibus[data_w*3 +:data_w] = c665obus[data_w*0 +:data_w];
assign c665ibus[temp_w*1 +:temp_w] = v334obus[temp_w*1 +:temp_w];
assign v334ibus[data_w*1 +:data_w] = c665obus[data_w*1 +:data_w];
assign c665ibus[temp_w*2 +:temp_w] = v871obus[temp_w*3 +:temp_w];
assign v871ibus[data_w*3 +:data_w] = c665obus[data_w*2 +:data_w];
assign c665ibus[temp_w*3 +:temp_w] = v971obus[temp_w*1 +:temp_w];
assign v971ibus[data_w*1 +:data_w] = c665obus[data_w*3 +:data_w];
assign c665ibus[temp_w*4 +:temp_w] = v1817obus[temp_w*1 +:temp_w];
assign v1817ibus[data_w*1 +:data_w] = c665obus[data_w*4 +:data_w];
assign c665ibus[temp_w*5 +:temp_w] = v1913obus[temp_w*0 +:temp_w];
assign v1913ibus[data_w*0 +:data_w] = c665obus[data_w*5 +:data_w];
assign c666ibus[temp_w*0 +:temp_w] = v281obus[temp_w*3 +:temp_w];
assign v281ibus[data_w*3 +:data_w] = c666obus[data_w*0 +:data_w];
assign c666ibus[temp_w*1 +:temp_w] = v335obus[temp_w*1 +:temp_w];
assign v335ibus[data_w*1 +:data_w] = c666obus[data_w*1 +:data_w];
assign c666ibus[temp_w*2 +:temp_w] = v872obus[temp_w*3 +:temp_w];
assign v872ibus[data_w*3 +:data_w] = c666obus[data_w*2 +:data_w];
assign c666ibus[temp_w*3 +:temp_w] = v972obus[temp_w*1 +:temp_w];
assign v972ibus[data_w*1 +:data_w] = c666obus[data_w*3 +:data_w];
assign c666ibus[temp_w*4 +:temp_w] = v1818obus[temp_w*1 +:temp_w];
assign v1818ibus[data_w*1 +:data_w] = c666obus[data_w*4 +:data_w];
assign c666ibus[temp_w*5 +:temp_w] = v1914obus[temp_w*0 +:temp_w];
assign v1914ibus[data_w*0 +:data_w] = c666obus[data_w*5 +:data_w];
assign c667ibus[temp_w*0 +:temp_w] = v282obus[temp_w*3 +:temp_w];
assign v282ibus[data_w*3 +:data_w] = c667obus[data_w*0 +:data_w];
assign c667ibus[temp_w*1 +:temp_w] = v336obus[temp_w*1 +:temp_w];
assign v336ibus[data_w*1 +:data_w] = c667obus[data_w*1 +:data_w];
assign c667ibus[temp_w*2 +:temp_w] = v873obus[temp_w*3 +:temp_w];
assign v873ibus[data_w*3 +:data_w] = c667obus[data_w*2 +:data_w];
assign c667ibus[temp_w*3 +:temp_w] = v973obus[temp_w*1 +:temp_w];
assign v973ibus[data_w*1 +:data_w] = c667obus[data_w*3 +:data_w];
assign c667ibus[temp_w*4 +:temp_w] = v1819obus[temp_w*1 +:temp_w];
assign v1819ibus[data_w*1 +:data_w] = c667obus[data_w*4 +:data_w];
assign c667ibus[temp_w*5 +:temp_w] = v1915obus[temp_w*0 +:temp_w];
assign v1915ibus[data_w*0 +:data_w] = c667obus[data_w*5 +:data_w];
assign c668ibus[temp_w*0 +:temp_w] = v283obus[temp_w*3 +:temp_w];
assign v283ibus[data_w*3 +:data_w] = c668obus[data_w*0 +:data_w];
assign c668ibus[temp_w*1 +:temp_w] = v337obus[temp_w*1 +:temp_w];
assign v337ibus[data_w*1 +:data_w] = c668obus[data_w*1 +:data_w];
assign c668ibus[temp_w*2 +:temp_w] = v874obus[temp_w*3 +:temp_w];
assign v874ibus[data_w*3 +:data_w] = c668obus[data_w*2 +:data_w];
assign c668ibus[temp_w*3 +:temp_w] = v974obus[temp_w*1 +:temp_w];
assign v974ibus[data_w*1 +:data_w] = c668obus[data_w*3 +:data_w];
assign c668ibus[temp_w*4 +:temp_w] = v1820obus[temp_w*1 +:temp_w];
assign v1820ibus[data_w*1 +:data_w] = c668obus[data_w*4 +:data_w];
assign c668ibus[temp_w*5 +:temp_w] = v1916obus[temp_w*0 +:temp_w];
assign v1916ibus[data_w*0 +:data_w] = c668obus[data_w*5 +:data_w];
assign c669ibus[temp_w*0 +:temp_w] = v284obus[temp_w*3 +:temp_w];
assign v284ibus[data_w*3 +:data_w] = c669obus[data_w*0 +:data_w];
assign c669ibus[temp_w*1 +:temp_w] = v338obus[temp_w*1 +:temp_w];
assign v338ibus[data_w*1 +:data_w] = c669obus[data_w*1 +:data_w];
assign c669ibus[temp_w*2 +:temp_w] = v875obus[temp_w*3 +:temp_w];
assign v875ibus[data_w*3 +:data_w] = c669obus[data_w*2 +:data_w];
assign c669ibus[temp_w*3 +:temp_w] = v975obus[temp_w*1 +:temp_w];
assign v975ibus[data_w*1 +:data_w] = c669obus[data_w*3 +:data_w];
assign c669ibus[temp_w*4 +:temp_w] = v1821obus[temp_w*1 +:temp_w];
assign v1821ibus[data_w*1 +:data_w] = c669obus[data_w*4 +:data_w];
assign c669ibus[temp_w*5 +:temp_w] = v1917obus[temp_w*0 +:temp_w];
assign v1917ibus[data_w*0 +:data_w] = c669obus[data_w*5 +:data_w];
assign c670ibus[temp_w*0 +:temp_w] = v285obus[temp_w*3 +:temp_w];
assign v285ibus[data_w*3 +:data_w] = c670obus[data_w*0 +:data_w];
assign c670ibus[temp_w*1 +:temp_w] = v339obus[temp_w*1 +:temp_w];
assign v339ibus[data_w*1 +:data_w] = c670obus[data_w*1 +:data_w];
assign c670ibus[temp_w*2 +:temp_w] = v876obus[temp_w*3 +:temp_w];
assign v876ibus[data_w*3 +:data_w] = c670obus[data_w*2 +:data_w];
assign c670ibus[temp_w*3 +:temp_w] = v976obus[temp_w*1 +:temp_w];
assign v976ibus[data_w*1 +:data_w] = c670obus[data_w*3 +:data_w];
assign c670ibus[temp_w*4 +:temp_w] = v1822obus[temp_w*1 +:temp_w];
assign v1822ibus[data_w*1 +:data_w] = c670obus[data_w*4 +:data_w];
assign c670ibus[temp_w*5 +:temp_w] = v1918obus[temp_w*0 +:temp_w];
assign v1918ibus[data_w*0 +:data_w] = c670obus[data_w*5 +:data_w];
assign c671ibus[temp_w*0 +:temp_w] = v286obus[temp_w*3 +:temp_w];
assign v286ibus[data_w*3 +:data_w] = c671obus[data_w*0 +:data_w];
assign c671ibus[temp_w*1 +:temp_w] = v340obus[temp_w*1 +:temp_w];
assign v340ibus[data_w*1 +:data_w] = c671obus[data_w*1 +:data_w];
assign c671ibus[temp_w*2 +:temp_w] = v877obus[temp_w*3 +:temp_w];
assign v877ibus[data_w*3 +:data_w] = c671obus[data_w*2 +:data_w];
assign c671ibus[temp_w*3 +:temp_w] = v977obus[temp_w*1 +:temp_w];
assign v977ibus[data_w*1 +:data_w] = c671obus[data_w*3 +:data_w];
assign c671ibus[temp_w*4 +:temp_w] = v1823obus[temp_w*1 +:temp_w];
assign v1823ibus[data_w*1 +:data_w] = c671obus[data_w*4 +:data_w];
assign c671ibus[temp_w*5 +:temp_w] = v1919obus[temp_w*0 +:temp_w];
assign v1919ibus[data_w*0 +:data_w] = c671obus[data_w*5 +:data_w];
assign c672ibus[temp_w*0 +:temp_w] = v107obus[temp_w*2 +:temp_w];
assign v107ibus[data_w*2 +:data_w] = c672obus[data_w*0 +:data_w];
assign c672ibus[temp_w*1 +:temp_w] = v265obus[temp_w*4 +:temp_w];
assign v265ibus[data_w*4 +:data_w] = c672obus[data_w*1 +:data_w];
assign c672ibus[temp_w*2 +:temp_w] = v578obus[temp_w*2 +:temp_w];
assign v578ibus[data_w*2 +:data_w] = c672obus[data_w*2 +:data_w];
assign c672ibus[temp_w*3 +:temp_w] = v911obus[temp_w*4 +:temp_w];
assign v911ibus[data_w*4 +:data_w] = c672obus[data_w*3 +:data_w];
assign c672ibus[temp_w*4 +:temp_w] = v1824obus[temp_w*1 +:temp_w];
assign v1824ibus[data_w*1 +:data_w] = c672obus[data_w*4 +:data_w];
assign c672ibus[temp_w*5 +:temp_w] = v1920obus[temp_w*0 +:temp_w];
assign v1920ibus[data_w*0 +:data_w] = c672obus[data_w*5 +:data_w];
assign c673ibus[temp_w*0 +:temp_w] = v108obus[temp_w*2 +:temp_w];
assign v108ibus[data_w*2 +:data_w] = c673obus[data_w*0 +:data_w];
assign c673ibus[temp_w*1 +:temp_w] = v266obus[temp_w*4 +:temp_w];
assign v266ibus[data_w*4 +:data_w] = c673obus[data_w*1 +:data_w];
assign c673ibus[temp_w*2 +:temp_w] = v579obus[temp_w*2 +:temp_w];
assign v579ibus[data_w*2 +:data_w] = c673obus[data_w*2 +:data_w];
assign c673ibus[temp_w*3 +:temp_w] = v912obus[temp_w*4 +:temp_w];
assign v912ibus[data_w*4 +:data_w] = c673obus[data_w*3 +:data_w];
assign c673ibus[temp_w*4 +:temp_w] = v1825obus[temp_w*1 +:temp_w];
assign v1825ibus[data_w*1 +:data_w] = c673obus[data_w*4 +:data_w];
assign c673ibus[temp_w*5 +:temp_w] = v1921obus[temp_w*0 +:temp_w];
assign v1921ibus[data_w*0 +:data_w] = c673obus[data_w*5 +:data_w];
assign c674ibus[temp_w*0 +:temp_w] = v109obus[temp_w*2 +:temp_w];
assign v109ibus[data_w*2 +:data_w] = c674obus[data_w*0 +:data_w];
assign c674ibus[temp_w*1 +:temp_w] = v267obus[temp_w*4 +:temp_w];
assign v267ibus[data_w*4 +:data_w] = c674obus[data_w*1 +:data_w];
assign c674ibus[temp_w*2 +:temp_w] = v580obus[temp_w*2 +:temp_w];
assign v580ibus[data_w*2 +:data_w] = c674obus[data_w*2 +:data_w];
assign c674ibus[temp_w*3 +:temp_w] = v913obus[temp_w*4 +:temp_w];
assign v913ibus[data_w*4 +:data_w] = c674obus[data_w*3 +:data_w];
assign c674ibus[temp_w*4 +:temp_w] = v1826obus[temp_w*1 +:temp_w];
assign v1826ibus[data_w*1 +:data_w] = c674obus[data_w*4 +:data_w];
assign c674ibus[temp_w*5 +:temp_w] = v1922obus[temp_w*0 +:temp_w];
assign v1922ibus[data_w*0 +:data_w] = c674obus[data_w*5 +:data_w];
assign c675ibus[temp_w*0 +:temp_w] = v110obus[temp_w*2 +:temp_w];
assign v110ibus[data_w*2 +:data_w] = c675obus[data_w*0 +:data_w];
assign c675ibus[temp_w*1 +:temp_w] = v268obus[temp_w*4 +:temp_w];
assign v268ibus[data_w*4 +:data_w] = c675obus[data_w*1 +:data_w];
assign c675ibus[temp_w*2 +:temp_w] = v581obus[temp_w*2 +:temp_w];
assign v581ibus[data_w*2 +:data_w] = c675obus[data_w*2 +:data_w];
assign c675ibus[temp_w*3 +:temp_w] = v914obus[temp_w*4 +:temp_w];
assign v914ibus[data_w*4 +:data_w] = c675obus[data_w*3 +:data_w];
assign c675ibus[temp_w*4 +:temp_w] = v1827obus[temp_w*1 +:temp_w];
assign v1827ibus[data_w*1 +:data_w] = c675obus[data_w*4 +:data_w];
assign c675ibus[temp_w*5 +:temp_w] = v1923obus[temp_w*0 +:temp_w];
assign v1923ibus[data_w*0 +:data_w] = c675obus[data_w*5 +:data_w];
assign c676ibus[temp_w*0 +:temp_w] = v111obus[temp_w*2 +:temp_w];
assign v111ibus[data_w*2 +:data_w] = c676obus[data_w*0 +:data_w];
assign c676ibus[temp_w*1 +:temp_w] = v269obus[temp_w*4 +:temp_w];
assign v269ibus[data_w*4 +:data_w] = c676obus[data_w*1 +:data_w];
assign c676ibus[temp_w*2 +:temp_w] = v582obus[temp_w*2 +:temp_w];
assign v582ibus[data_w*2 +:data_w] = c676obus[data_w*2 +:data_w];
assign c676ibus[temp_w*3 +:temp_w] = v915obus[temp_w*4 +:temp_w];
assign v915ibus[data_w*4 +:data_w] = c676obus[data_w*3 +:data_w];
assign c676ibus[temp_w*4 +:temp_w] = v1828obus[temp_w*1 +:temp_w];
assign v1828ibus[data_w*1 +:data_w] = c676obus[data_w*4 +:data_w];
assign c676ibus[temp_w*5 +:temp_w] = v1924obus[temp_w*0 +:temp_w];
assign v1924ibus[data_w*0 +:data_w] = c676obus[data_w*5 +:data_w];
assign c677ibus[temp_w*0 +:temp_w] = v112obus[temp_w*2 +:temp_w];
assign v112ibus[data_w*2 +:data_w] = c677obus[data_w*0 +:data_w];
assign c677ibus[temp_w*1 +:temp_w] = v270obus[temp_w*4 +:temp_w];
assign v270ibus[data_w*4 +:data_w] = c677obus[data_w*1 +:data_w];
assign c677ibus[temp_w*2 +:temp_w] = v583obus[temp_w*2 +:temp_w];
assign v583ibus[data_w*2 +:data_w] = c677obus[data_w*2 +:data_w];
assign c677ibus[temp_w*3 +:temp_w] = v916obus[temp_w*4 +:temp_w];
assign v916ibus[data_w*4 +:data_w] = c677obus[data_w*3 +:data_w];
assign c677ibus[temp_w*4 +:temp_w] = v1829obus[temp_w*1 +:temp_w];
assign v1829ibus[data_w*1 +:data_w] = c677obus[data_w*4 +:data_w];
assign c677ibus[temp_w*5 +:temp_w] = v1925obus[temp_w*0 +:temp_w];
assign v1925ibus[data_w*0 +:data_w] = c677obus[data_w*5 +:data_w];
assign c678ibus[temp_w*0 +:temp_w] = v113obus[temp_w*2 +:temp_w];
assign v113ibus[data_w*2 +:data_w] = c678obus[data_w*0 +:data_w];
assign c678ibus[temp_w*1 +:temp_w] = v271obus[temp_w*4 +:temp_w];
assign v271ibus[data_w*4 +:data_w] = c678obus[data_w*1 +:data_w];
assign c678ibus[temp_w*2 +:temp_w] = v584obus[temp_w*2 +:temp_w];
assign v584ibus[data_w*2 +:data_w] = c678obus[data_w*2 +:data_w];
assign c678ibus[temp_w*3 +:temp_w] = v917obus[temp_w*4 +:temp_w];
assign v917ibus[data_w*4 +:data_w] = c678obus[data_w*3 +:data_w];
assign c678ibus[temp_w*4 +:temp_w] = v1830obus[temp_w*1 +:temp_w];
assign v1830ibus[data_w*1 +:data_w] = c678obus[data_w*4 +:data_w];
assign c678ibus[temp_w*5 +:temp_w] = v1926obus[temp_w*0 +:temp_w];
assign v1926ibus[data_w*0 +:data_w] = c678obus[data_w*5 +:data_w];
assign c679ibus[temp_w*0 +:temp_w] = v114obus[temp_w*2 +:temp_w];
assign v114ibus[data_w*2 +:data_w] = c679obus[data_w*0 +:data_w];
assign c679ibus[temp_w*1 +:temp_w] = v272obus[temp_w*4 +:temp_w];
assign v272ibus[data_w*4 +:data_w] = c679obus[data_w*1 +:data_w];
assign c679ibus[temp_w*2 +:temp_w] = v585obus[temp_w*2 +:temp_w];
assign v585ibus[data_w*2 +:data_w] = c679obus[data_w*2 +:data_w];
assign c679ibus[temp_w*3 +:temp_w] = v918obus[temp_w*4 +:temp_w];
assign v918ibus[data_w*4 +:data_w] = c679obus[data_w*3 +:data_w];
assign c679ibus[temp_w*4 +:temp_w] = v1831obus[temp_w*1 +:temp_w];
assign v1831ibus[data_w*1 +:data_w] = c679obus[data_w*4 +:data_w];
assign c679ibus[temp_w*5 +:temp_w] = v1927obus[temp_w*0 +:temp_w];
assign v1927ibus[data_w*0 +:data_w] = c679obus[data_w*5 +:data_w];
assign c680ibus[temp_w*0 +:temp_w] = v115obus[temp_w*2 +:temp_w];
assign v115ibus[data_w*2 +:data_w] = c680obus[data_w*0 +:data_w];
assign c680ibus[temp_w*1 +:temp_w] = v273obus[temp_w*4 +:temp_w];
assign v273ibus[data_w*4 +:data_w] = c680obus[data_w*1 +:data_w];
assign c680ibus[temp_w*2 +:temp_w] = v586obus[temp_w*2 +:temp_w];
assign v586ibus[data_w*2 +:data_w] = c680obus[data_w*2 +:data_w];
assign c680ibus[temp_w*3 +:temp_w] = v919obus[temp_w*4 +:temp_w];
assign v919ibus[data_w*4 +:data_w] = c680obus[data_w*3 +:data_w];
assign c680ibus[temp_w*4 +:temp_w] = v1832obus[temp_w*1 +:temp_w];
assign v1832ibus[data_w*1 +:data_w] = c680obus[data_w*4 +:data_w];
assign c680ibus[temp_w*5 +:temp_w] = v1928obus[temp_w*0 +:temp_w];
assign v1928ibus[data_w*0 +:data_w] = c680obus[data_w*5 +:data_w];
assign c681ibus[temp_w*0 +:temp_w] = v116obus[temp_w*2 +:temp_w];
assign v116ibus[data_w*2 +:data_w] = c681obus[data_w*0 +:data_w];
assign c681ibus[temp_w*1 +:temp_w] = v274obus[temp_w*4 +:temp_w];
assign v274ibus[data_w*4 +:data_w] = c681obus[data_w*1 +:data_w];
assign c681ibus[temp_w*2 +:temp_w] = v587obus[temp_w*2 +:temp_w];
assign v587ibus[data_w*2 +:data_w] = c681obus[data_w*2 +:data_w];
assign c681ibus[temp_w*3 +:temp_w] = v920obus[temp_w*4 +:temp_w];
assign v920ibus[data_w*4 +:data_w] = c681obus[data_w*3 +:data_w];
assign c681ibus[temp_w*4 +:temp_w] = v1833obus[temp_w*1 +:temp_w];
assign v1833ibus[data_w*1 +:data_w] = c681obus[data_w*4 +:data_w];
assign c681ibus[temp_w*5 +:temp_w] = v1929obus[temp_w*0 +:temp_w];
assign v1929ibus[data_w*0 +:data_w] = c681obus[data_w*5 +:data_w];
assign c682ibus[temp_w*0 +:temp_w] = v117obus[temp_w*2 +:temp_w];
assign v117ibus[data_w*2 +:data_w] = c682obus[data_w*0 +:data_w];
assign c682ibus[temp_w*1 +:temp_w] = v275obus[temp_w*4 +:temp_w];
assign v275ibus[data_w*4 +:data_w] = c682obus[data_w*1 +:data_w];
assign c682ibus[temp_w*2 +:temp_w] = v588obus[temp_w*2 +:temp_w];
assign v588ibus[data_w*2 +:data_w] = c682obus[data_w*2 +:data_w];
assign c682ibus[temp_w*3 +:temp_w] = v921obus[temp_w*4 +:temp_w];
assign v921ibus[data_w*4 +:data_w] = c682obus[data_w*3 +:data_w];
assign c682ibus[temp_w*4 +:temp_w] = v1834obus[temp_w*1 +:temp_w];
assign v1834ibus[data_w*1 +:data_w] = c682obus[data_w*4 +:data_w];
assign c682ibus[temp_w*5 +:temp_w] = v1930obus[temp_w*0 +:temp_w];
assign v1930ibus[data_w*0 +:data_w] = c682obus[data_w*5 +:data_w];
assign c683ibus[temp_w*0 +:temp_w] = v118obus[temp_w*2 +:temp_w];
assign v118ibus[data_w*2 +:data_w] = c683obus[data_w*0 +:data_w];
assign c683ibus[temp_w*1 +:temp_w] = v276obus[temp_w*4 +:temp_w];
assign v276ibus[data_w*4 +:data_w] = c683obus[data_w*1 +:data_w];
assign c683ibus[temp_w*2 +:temp_w] = v589obus[temp_w*2 +:temp_w];
assign v589ibus[data_w*2 +:data_w] = c683obus[data_w*2 +:data_w];
assign c683ibus[temp_w*3 +:temp_w] = v922obus[temp_w*4 +:temp_w];
assign v922ibus[data_w*4 +:data_w] = c683obus[data_w*3 +:data_w];
assign c683ibus[temp_w*4 +:temp_w] = v1835obus[temp_w*1 +:temp_w];
assign v1835ibus[data_w*1 +:data_w] = c683obus[data_w*4 +:data_w];
assign c683ibus[temp_w*5 +:temp_w] = v1931obus[temp_w*0 +:temp_w];
assign v1931ibus[data_w*0 +:data_w] = c683obus[data_w*5 +:data_w];
assign c684ibus[temp_w*0 +:temp_w] = v119obus[temp_w*2 +:temp_w];
assign v119ibus[data_w*2 +:data_w] = c684obus[data_w*0 +:data_w];
assign c684ibus[temp_w*1 +:temp_w] = v277obus[temp_w*4 +:temp_w];
assign v277ibus[data_w*4 +:data_w] = c684obus[data_w*1 +:data_w];
assign c684ibus[temp_w*2 +:temp_w] = v590obus[temp_w*2 +:temp_w];
assign v590ibus[data_w*2 +:data_w] = c684obus[data_w*2 +:data_w];
assign c684ibus[temp_w*3 +:temp_w] = v923obus[temp_w*4 +:temp_w];
assign v923ibus[data_w*4 +:data_w] = c684obus[data_w*3 +:data_w];
assign c684ibus[temp_w*4 +:temp_w] = v1836obus[temp_w*1 +:temp_w];
assign v1836ibus[data_w*1 +:data_w] = c684obus[data_w*4 +:data_w];
assign c684ibus[temp_w*5 +:temp_w] = v1932obus[temp_w*0 +:temp_w];
assign v1932ibus[data_w*0 +:data_w] = c684obus[data_w*5 +:data_w];
assign c685ibus[temp_w*0 +:temp_w] = v120obus[temp_w*2 +:temp_w];
assign v120ibus[data_w*2 +:data_w] = c685obus[data_w*0 +:data_w];
assign c685ibus[temp_w*1 +:temp_w] = v278obus[temp_w*4 +:temp_w];
assign v278ibus[data_w*4 +:data_w] = c685obus[data_w*1 +:data_w];
assign c685ibus[temp_w*2 +:temp_w] = v591obus[temp_w*2 +:temp_w];
assign v591ibus[data_w*2 +:data_w] = c685obus[data_w*2 +:data_w];
assign c685ibus[temp_w*3 +:temp_w] = v924obus[temp_w*4 +:temp_w];
assign v924ibus[data_w*4 +:data_w] = c685obus[data_w*3 +:data_w];
assign c685ibus[temp_w*4 +:temp_w] = v1837obus[temp_w*1 +:temp_w];
assign v1837ibus[data_w*1 +:data_w] = c685obus[data_w*4 +:data_w];
assign c685ibus[temp_w*5 +:temp_w] = v1933obus[temp_w*0 +:temp_w];
assign v1933ibus[data_w*0 +:data_w] = c685obus[data_w*5 +:data_w];
assign c686ibus[temp_w*0 +:temp_w] = v121obus[temp_w*2 +:temp_w];
assign v121ibus[data_w*2 +:data_w] = c686obus[data_w*0 +:data_w];
assign c686ibus[temp_w*1 +:temp_w] = v279obus[temp_w*4 +:temp_w];
assign v279ibus[data_w*4 +:data_w] = c686obus[data_w*1 +:data_w];
assign c686ibus[temp_w*2 +:temp_w] = v592obus[temp_w*2 +:temp_w];
assign v592ibus[data_w*2 +:data_w] = c686obus[data_w*2 +:data_w];
assign c686ibus[temp_w*3 +:temp_w] = v925obus[temp_w*4 +:temp_w];
assign v925ibus[data_w*4 +:data_w] = c686obus[data_w*3 +:data_w];
assign c686ibus[temp_w*4 +:temp_w] = v1838obus[temp_w*1 +:temp_w];
assign v1838ibus[data_w*1 +:data_w] = c686obus[data_w*4 +:data_w];
assign c686ibus[temp_w*5 +:temp_w] = v1934obus[temp_w*0 +:temp_w];
assign v1934ibus[data_w*0 +:data_w] = c686obus[data_w*5 +:data_w];
assign c687ibus[temp_w*0 +:temp_w] = v122obus[temp_w*2 +:temp_w];
assign v122ibus[data_w*2 +:data_w] = c687obus[data_w*0 +:data_w];
assign c687ibus[temp_w*1 +:temp_w] = v280obus[temp_w*4 +:temp_w];
assign v280ibus[data_w*4 +:data_w] = c687obus[data_w*1 +:data_w];
assign c687ibus[temp_w*2 +:temp_w] = v593obus[temp_w*2 +:temp_w];
assign v593ibus[data_w*2 +:data_w] = c687obus[data_w*2 +:data_w];
assign c687ibus[temp_w*3 +:temp_w] = v926obus[temp_w*4 +:temp_w];
assign v926ibus[data_w*4 +:data_w] = c687obus[data_w*3 +:data_w];
assign c687ibus[temp_w*4 +:temp_w] = v1839obus[temp_w*1 +:temp_w];
assign v1839ibus[data_w*1 +:data_w] = c687obus[data_w*4 +:data_w];
assign c687ibus[temp_w*5 +:temp_w] = v1935obus[temp_w*0 +:temp_w];
assign v1935ibus[data_w*0 +:data_w] = c687obus[data_w*5 +:data_w];
assign c688ibus[temp_w*0 +:temp_w] = v123obus[temp_w*2 +:temp_w];
assign v123ibus[data_w*2 +:data_w] = c688obus[data_w*0 +:data_w];
assign c688ibus[temp_w*1 +:temp_w] = v281obus[temp_w*4 +:temp_w];
assign v281ibus[data_w*4 +:data_w] = c688obus[data_w*1 +:data_w];
assign c688ibus[temp_w*2 +:temp_w] = v594obus[temp_w*2 +:temp_w];
assign v594ibus[data_w*2 +:data_w] = c688obus[data_w*2 +:data_w];
assign c688ibus[temp_w*3 +:temp_w] = v927obus[temp_w*4 +:temp_w];
assign v927ibus[data_w*4 +:data_w] = c688obus[data_w*3 +:data_w];
assign c688ibus[temp_w*4 +:temp_w] = v1840obus[temp_w*1 +:temp_w];
assign v1840ibus[data_w*1 +:data_w] = c688obus[data_w*4 +:data_w];
assign c688ibus[temp_w*5 +:temp_w] = v1936obus[temp_w*0 +:temp_w];
assign v1936ibus[data_w*0 +:data_w] = c688obus[data_w*5 +:data_w];
assign c689ibus[temp_w*0 +:temp_w] = v124obus[temp_w*2 +:temp_w];
assign v124ibus[data_w*2 +:data_w] = c689obus[data_w*0 +:data_w];
assign c689ibus[temp_w*1 +:temp_w] = v282obus[temp_w*4 +:temp_w];
assign v282ibus[data_w*4 +:data_w] = c689obus[data_w*1 +:data_w];
assign c689ibus[temp_w*2 +:temp_w] = v595obus[temp_w*2 +:temp_w];
assign v595ibus[data_w*2 +:data_w] = c689obus[data_w*2 +:data_w];
assign c689ibus[temp_w*3 +:temp_w] = v928obus[temp_w*4 +:temp_w];
assign v928ibus[data_w*4 +:data_w] = c689obus[data_w*3 +:data_w];
assign c689ibus[temp_w*4 +:temp_w] = v1841obus[temp_w*1 +:temp_w];
assign v1841ibus[data_w*1 +:data_w] = c689obus[data_w*4 +:data_w];
assign c689ibus[temp_w*5 +:temp_w] = v1937obus[temp_w*0 +:temp_w];
assign v1937ibus[data_w*0 +:data_w] = c689obus[data_w*5 +:data_w];
assign c690ibus[temp_w*0 +:temp_w] = v125obus[temp_w*2 +:temp_w];
assign v125ibus[data_w*2 +:data_w] = c690obus[data_w*0 +:data_w];
assign c690ibus[temp_w*1 +:temp_w] = v283obus[temp_w*4 +:temp_w];
assign v283ibus[data_w*4 +:data_w] = c690obus[data_w*1 +:data_w];
assign c690ibus[temp_w*2 +:temp_w] = v596obus[temp_w*2 +:temp_w];
assign v596ibus[data_w*2 +:data_w] = c690obus[data_w*2 +:data_w];
assign c690ibus[temp_w*3 +:temp_w] = v929obus[temp_w*4 +:temp_w];
assign v929ibus[data_w*4 +:data_w] = c690obus[data_w*3 +:data_w];
assign c690ibus[temp_w*4 +:temp_w] = v1842obus[temp_w*1 +:temp_w];
assign v1842ibus[data_w*1 +:data_w] = c690obus[data_w*4 +:data_w];
assign c690ibus[temp_w*5 +:temp_w] = v1938obus[temp_w*0 +:temp_w];
assign v1938ibus[data_w*0 +:data_w] = c690obus[data_w*5 +:data_w];
assign c691ibus[temp_w*0 +:temp_w] = v126obus[temp_w*2 +:temp_w];
assign v126ibus[data_w*2 +:data_w] = c691obus[data_w*0 +:data_w];
assign c691ibus[temp_w*1 +:temp_w] = v284obus[temp_w*4 +:temp_w];
assign v284ibus[data_w*4 +:data_w] = c691obus[data_w*1 +:data_w];
assign c691ibus[temp_w*2 +:temp_w] = v597obus[temp_w*2 +:temp_w];
assign v597ibus[data_w*2 +:data_w] = c691obus[data_w*2 +:data_w];
assign c691ibus[temp_w*3 +:temp_w] = v930obus[temp_w*4 +:temp_w];
assign v930ibus[data_w*4 +:data_w] = c691obus[data_w*3 +:data_w];
assign c691ibus[temp_w*4 +:temp_w] = v1843obus[temp_w*1 +:temp_w];
assign v1843ibus[data_w*1 +:data_w] = c691obus[data_w*4 +:data_w];
assign c691ibus[temp_w*5 +:temp_w] = v1939obus[temp_w*0 +:temp_w];
assign v1939ibus[data_w*0 +:data_w] = c691obus[data_w*5 +:data_w];
assign c692ibus[temp_w*0 +:temp_w] = v127obus[temp_w*2 +:temp_w];
assign v127ibus[data_w*2 +:data_w] = c692obus[data_w*0 +:data_w];
assign c692ibus[temp_w*1 +:temp_w] = v285obus[temp_w*4 +:temp_w];
assign v285ibus[data_w*4 +:data_w] = c692obus[data_w*1 +:data_w];
assign c692ibus[temp_w*2 +:temp_w] = v598obus[temp_w*2 +:temp_w];
assign v598ibus[data_w*2 +:data_w] = c692obus[data_w*2 +:data_w];
assign c692ibus[temp_w*3 +:temp_w] = v931obus[temp_w*4 +:temp_w];
assign v931ibus[data_w*4 +:data_w] = c692obus[data_w*3 +:data_w];
assign c692ibus[temp_w*4 +:temp_w] = v1844obus[temp_w*1 +:temp_w];
assign v1844ibus[data_w*1 +:data_w] = c692obus[data_w*4 +:data_w];
assign c692ibus[temp_w*5 +:temp_w] = v1940obus[temp_w*0 +:temp_w];
assign v1940ibus[data_w*0 +:data_w] = c692obus[data_w*5 +:data_w];
assign c693ibus[temp_w*0 +:temp_w] = v128obus[temp_w*2 +:temp_w];
assign v128ibus[data_w*2 +:data_w] = c693obus[data_w*0 +:data_w];
assign c693ibus[temp_w*1 +:temp_w] = v286obus[temp_w*4 +:temp_w];
assign v286ibus[data_w*4 +:data_w] = c693obus[data_w*1 +:data_w];
assign c693ibus[temp_w*2 +:temp_w] = v599obus[temp_w*2 +:temp_w];
assign v599ibus[data_w*2 +:data_w] = c693obus[data_w*2 +:data_w];
assign c693ibus[temp_w*3 +:temp_w] = v932obus[temp_w*4 +:temp_w];
assign v932ibus[data_w*4 +:data_w] = c693obus[data_w*3 +:data_w];
assign c693ibus[temp_w*4 +:temp_w] = v1845obus[temp_w*1 +:temp_w];
assign v1845ibus[data_w*1 +:data_w] = c693obus[data_w*4 +:data_w];
assign c693ibus[temp_w*5 +:temp_w] = v1941obus[temp_w*0 +:temp_w];
assign v1941ibus[data_w*0 +:data_w] = c693obus[data_w*5 +:data_w];
assign c694ibus[temp_w*0 +:temp_w] = v129obus[temp_w*2 +:temp_w];
assign v129ibus[data_w*2 +:data_w] = c694obus[data_w*0 +:data_w];
assign c694ibus[temp_w*1 +:temp_w] = v287obus[temp_w*4 +:temp_w];
assign v287ibus[data_w*4 +:data_w] = c694obus[data_w*1 +:data_w];
assign c694ibus[temp_w*2 +:temp_w] = v600obus[temp_w*2 +:temp_w];
assign v600ibus[data_w*2 +:data_w] = c694obus[data_w*2 +:data_w];
assign c694ibus[temp_w*3 +:temp_w] = v933obus[temp_w*4 +:temp_w];
assign v933ibus[data_w*4 +:data_w] = c694obus[data_w*3 +:data_w];
assign c694ibus[temp_w*4 +:temp_w] = v1846obus[temp_w*1 +:temp_w];
assign v1846ibus[data_w*1 +:data_w] = c694obus[data_w*4 +:data_w];
assign c694ibus[temp_w*5 +:temp_w] = v1942obus[temp_w*0 +:temp_w];
assign v1942ibus[data_w*0 +:data_w] = c694obus[data_w*5 +:data_w];
assign c695ibus[temp_w*0 +:temp_w] = v130obus[temp_w*2 +:temp_w];
assign v130ibus[data_w*2 +:data_w] = c695obus[data_w*0 +:data_w];
assign c695ibus[temp_w*1 +:temp_w] = v192obus[temp_w*4 +:temp_w];
assign v192ibus[data_w*4 +:data_w] = c695obus[data_w*1 +:data_w];
assign c695ibus[temp_w*2 +:temp_w] = v601obus[temp_w*2 +:temp_w];
assign v601ibus[data_w*2 +:data_w] = c695obus[data_w*2 +:data_w];
assign c695ibus[temp_w*3 +:temp_w] = v934obus[temp_w*4 +:temp_w];
assign v934ibus[data_w*4 +:data_w] = c695obus[data_w*3 +:data_w];
assign c695ibus[temp_w*4 +:temp_w] = v1847obus[temp_w*1 +:temp_w];
assign v1847ibus[data_w*1 +:data_w] = c695obus[data_w*4 +:data_w];
assign c695ibus[temp_w*5 +:temp_w] = v1943obus[temp_w*0 +:temp_w];
assign v1943ibus[data_w*0 +:data_w] = c695obus[data_w*5 +:data_w];
assign c696ibus[temp_w*0 +:temp_w] = v131obus[temp_w*2 +:temp_w];
assign v131ibus[data_w*2 +:data_w] = c696obus[data_w*0 +:data_w];
assign c696ibus[temp_w*1 +:temp_w] = v193obus[temp_w*4 +:temp_w];
assign v193ibus[data_w*4 +:data_w] = c696obus[data_w*1 +:data_w];
assign c696ibus[temp_w*2 +:temp_w] = v602obus[temp_w*2 +:temp_w];
assign v602ibus[data_w*2 +:data_w] = c696obus[data_w*2 +:data_w];
assign c696ibus[temp_w*3 +:temp_w] = v935obus[temp_w*4 +:temp_w];
assign v935ibus[data_w*4 +:data_w] = c696obus[data_w*3 +:data_w];
assign c696ibus[temp_w*4 +:temp_w] = v1848obus[temp_w*1 +:temp_w];
assign v1848ibus[data_w*1 +:data_w] = c696obus[data_w*4 +:data_w];
assign c696ibus[temp_w*5 +:temp_w] = v1944obus[temp_w*0 +:temp_w];
assign v1944ibus[data_w*0 +:data_w] = c696obus[data_w*5 +:data_w];
assign c697ibus[temp_w*0 +:temp_w] = v132obus[temp_w*2 +:temp_w];
assign v132ibus[data_w*2 +:data_w] = c697obus[data_w*0 +:data_w];
assign c697ibus[temp_w*1 +:temp_w] = v194obus[temp_w*4 +:temp_w];
assign v194ibus[data_w*4 +:data_w] = c697obus[data_w*1 +:data_w];
assign c697ibus[temp_w*2 +:temp_w] = v603obus[temp_w*2 +:temp_w];
assign v603ibus[data_w*2 +:data_w] = c697obus[data_w*2 +:data_w];
assign c697ibus[temp_w*3 +:temp_w] = v936obus[temp_w*4 +:temp_w];
assign v936ibus[data_w*4 +:data_w] = c697obus[data_w*3 +:data_w];
assign c697ibus[temp_w*4 +:temp_w] = v1849obus[temp_w*1 +:temp_w];
assign v1849ibus[data_w*1 +:data_w] = c697obus[data_w*4 +:data_w];
assign c697ibus[temp_w*5 +:temp_w] = v1945obus[temp_w*0 +:temp_w];
assign v1945ibus[data_w*0 +:data_w] = c697obus[data_w*5 +:data_w];
assign c698ibus[temp_w*0 +:temp_w] = v133obus[temp_w*2 +:temp_w];
assign v133ibus[data_w*2 +:data_w] = c698obus[data_w*0 +:data_w];
assign c698ibus[temp_w*1 +:temp_w] = v195obus[temp_w*4 +:temp_w];
assign v195ibus[data_w*4 +:data_w] = c698obus[data_w*1 +:data_w];
assign c698ibus[temp_w*2 +:temp_w] = v604obus[temp_w*2 +:temp_w];
assign v604ibus[data_w*2 +:data_w] = c698obus[data_w*2 +:data_w];
assign c698ibus[temp_w*3 +:temp_w] = v937obus[temp_w*4 +:temp_w];
assign v937ibus[data_w*4 +:data_w] = c698obus[data_w*3 +:data_w];
assign c698ibus[temp_w*4 +:temp_w] = v1850obus[temp_w*1 +:temp_w];
assign v1850ibus[data_w*1 +:data_w] = c698obus[data_w*4 +:data_w];
assign c698ibus[temp_w*5 +:temp_w] = v1946obus[temp_w*0 +:temp_w];
assign v1946ibus[data_w*0 +:data_w] = c698obus[data_w*5 +:data_w];
assign c699ibus[temp_w*0 +:temp_w] = v134obus[temp_w*2 +:temp_w];
assign v134ibus[data_w*2 +:data_w] = c699obus[data_w*0 +:data_w];
assign c699ibus[temp_w*1 +:temp_w] = v196obus[temp_w*4 +:temp_w];
assign v196ibus[data_w*4 +:data_w] = c699obus[data_w*1 +:data_w];
assign c699ibus[temp_w*2 +:temp_w] = v605obus[temp_w*2 +:temp_w];
assign v605ibus[data_w*2 +:data_w] = c699obus[data_w*2 +:data_w];
assign c699ibus[temp_w*3 +:temp_w] = v938obus[temp_w*4 +:temp_w];
assign v938ibus[data_w*4 +:data_w] = c699obus[data_w*3 +:data_w];
assign c699ibus[temp_w*4 +:temp_w] = v1851obus[temp_w*1 +:temp_w];
assign v1851ibus[data_w*1 +:data_w] = c699obus[data_w*4 +:data_w];
assign c699ibus[temp_w*5 +:temp_w] = v1947obus[temp_w*0 +:temp_w];
assign v1947ibus[data_w*0 +:data_w] = c699obus[data_w*5 +:data_w];
assign c700ibus[temp_w*0 +:temp_w] = v135obus[temp_w*2 +:temp_w];
assign v135ibus[data_w*2 +:data_w] = c700obus[data_w*0 +:data_w];
assign c700ibus[temp_w*1 +:temp_w] = v197obus[temp_w*4 +:temp_w];
assign v197ibus[data_w*4 +:data_w] = c700obus[data_w*1 +:data_w];
assign c700ibus[temp_w*2 +:temp_w] = v606obus[temp_w*2 +:temp_w];
assign v606ibus[data_w*2 +:data_w] = c700obus[data_w*2 +:data_w];
assign c700ibus[temp_w*3 +:temp_w] = v939obus[temp_w*4 +:temp_w];
assign v939ibus[data_w*4 +:data_w] = c700obus[data_w*3 +:data_w];
assign c700ibus[temp_w*4 +:temp_w] = v1852obus[temp_w*1 +:temp_w];
assign v1852ibus[data_w*1 +:data_w] = c700obus[data_w*4 +:data_w];
assign c700ibus[temp_w*5 +:temp_w] = v1948obus[temp_w*0 +:temp_w];
assign v1948ibus[data_w*0 +:data_w] = c700obus[data_w*5 +:data_w];
assign c701ibus[temp_w*0 +:temp_w] = v136obus[temp_w*2 +:temp_w];
assign v136ibus[data_w*2 +:data_w] = c701obus[data_w*0 +:data_w];
assign c701ibus[temp_w*1 +:temp_w] = v198obus[temp_w*4 +:temp_w];
assign v198ibus[data_w*4 +:data_w] = c701obus[data_w*1 +:data_w];
assign c701ibus[temp_w*2 +:temp_w] = v607obus[temp_w*2 +:temp_w];
assign v607ibus[data_w*2 +:data_w] = c701obus[data_w*2 +:data_w];
assign c701ibus[temp_w*3 +:temp_w] = v940obus[temp_w*4 +:temp_w];
assign v940ibus[data_w*4 +:data_w] = c701obus[data_w*3 +:data_w];
assign c701ibus[temp_w*4 +:temp_w] = v1853obus[temp_w*1 +:temp_w];
assign v1853ibus[data_w*1 +:data_w] = c701obus[data_w*4 +:data_w];
assign c701ibus[temp_w*5 +:temp_w] = v1949obus[temp_w*0 +:temp_w];
assign v1949ibus[data_w*0 +:data_w] = c701obus[data_w*5 +:data_w];
assign c702ibus[temp_w*0 +:temp_w] = v137obus[temp_w*2 +:temp_w];
assign v137ibus[data_w*2 +:data_w] = c702obus[data_w*0 +:data_w];
assign c702ibus[temp_w*1 +:temp_w] = v199obus[temp_w*4 +:temp_w];
assign v199ibus[data_w*4 +:data_w] = c702obus[data_w*1 +:data_w];
assign c702ibus[temp_w*2 +:temp_w] = v608obus[temp_w*2 +:temp_w];
assign v608ibus[data_w*2 +:data_w] = c702obus[data_w*2 +:data_w];
assign c702ibus[temp_w*3 +:temp_w] = v941obus[temp_w*4 +:temp_w];
assign v941ibus[data_w*4 +:data_w] = c702obus[data_w*3 +:data_w];
assign c702ibus[temp_w*4 +:temp_w] = v1854obus[temp_w*1 +:temp_w];
assign v1854ibus[data_w*1 +:data_w] = c702obus[data_w*4 +:data_w];
assign c702ibus[temp_w*5 +:temp_w] = v1950obus[temp_w*0 +:temp_w];
assign v1950ibus[data_w*0 +:data_w] = c702obus[data_w*5 +:data_w];
assign c703ibus[temp_w*0 +:temp_w] = v138obus[temp_w*2 +:temp_w];
assign v138ibus[data_w*2 +:data_w] = c703obus[data_w*0 +:data_w];
assign c703ibus[temp_w*1 +:temp_w] = v200obus[temp_w*4 +:temp_w];
assign v200ibus[data_w*4 +:data_w] = c703obus[data_w*1 +:data_w];
assign c703ibus[temp_w*2 +:temp_w] = v609obus[temp_w*2 +:temp_w];
assign v609ibus[data_w*2 +:data_w] = c703obus[data_w*2 +:data_w];
assign c703ibus[temp_w*3 +:temp_w] = v942obus[temp_w*4 +:temp_w];
assign v942ibus[data_w*4 +:data_w] = c703obus[data_w*3 +:data_w];
assign c703ibus[temp_w*4 +:temp_w] = v1855obus[temp_w*1 +:temp_w];
assign v1855ibus[data_w*1 +:data_w] = c703obus[data_w*4 +:data_w];
assign c703ibus[temp_w*5 +:temp_w] = v1951obus[temp_w*0 +:temp_w];
assign v1951ibus[data_w*0 +:data_w] = c703obus[data_w*5 +:data_w];
assign c704ibus[temp_w*0 +:temp_w] = v139obus[temp_w*2 +:temp_w];
assign v139ibus[data_w*2 +:data_w] = c704obus[data_w*0 +:data_w];
assign c704ibus[temp_w*1 +:temp_w] = v201obus[temp_w*4 +:temp_w];
assign v201ibus[data_w*4 +:data_w] = c704obus[data_w*1 +:data_w];
assign c704ibus[temp_w*2 +:temp_w] = v610obus[temp_w*2 +:temp_w];
assign v610ibus[data_w*2 +:data_w] = c704obus[data_w*2 +:data_w];
assign c704ibus[temp_w*3 +:temp_w] = v943obus[temp_w*4 +:temp_w];
assign v943ibus[data_w*4 +:data_w] = c704obus[data_w*3 +:data_w];
assign c704ibus[temp_w*4 +:temp_w] = v1856obus[temp_w*1 +:temp_w];
assign v1856ibus[data_w*1 +:data_w] = c704obus[data_w*4 +:data_w];
assign c704ibus[temp_w*5 +:temp_w] = v1952obus[temp_w*0 +:temp_w];
assign v1952ibus[data_w*0 +:data_w] = c704obus[data_w*5 +:data_w];
assign c705ibus[temp_w*0 +:temp_w] = v140obus[temp_w*2 +:temp_w];
assign v140ibus[data_w*2 +:data_w] = c705obus[data_w*0 +:data_w];
assign c705ibus[temp_w*1 +:temp_w] = v202obus[temp_w*4 +:temp_w];
assign v202ibus[data_w*4 +:data_w] = c705obus[data_w*1 +:data_w];
assign c705ibus[temp_w*2 +:temp_w] = v611obus[temp_w*2 +:temp_w];
assign v611ibus[data_w*2 +:data_w] = c705obus[data_w*2 +:data_w];
assign c705ibus[temp_w*3 +:temp_w] = v944obus[temp_w*4 +:temp_w];
assign v944ibus[data_w*4 +:data_w] = c705obus[data_w*3 +:data_w];
assign c705ibus[temp_w*4 +:temp_w] = v1857obus[temp_w*1 +:temp_w];
assign v1857ibus[data_w*1 +:data_w] = c705obus[data_w*4 +:data_w];
assign c705ibus[temp_w*5 +:temp_w] = v1953obus[temp_w*0 +:temp_w];
assign v1953ibus[data_w*0 +:data_w] = c705obus[data_w*5 +:data_w];
assign c706ibus[temp_w*0 +:temp_w] = v141obus[temp_w*2 +:temp_w];
assign v141ibus[data_w*2 +:data_w] = c706obus[data_w*0 +:data_w];
assign c706ibus[temp_w*1 +:temp_w] = v203obus[temp_w*4 +:temp_w];
assign v203ibus[data_w*4 +:data_w] = c706obus[data_w*1 +:data_w];
assign c706ibus[temp_w*2 +:temp_w] = v612obus[temp_w*2 +:temp_w];
assign v612ibus[data_w*2 +:data_w] = c706obus[data_w*2 +:data_w];
assign c706ibus[temp_w*3 +:temp_w] = v945obus[temp_w*4 +:temp_w];
assign v945ibus[data_w*4 +:data_w] = c706obus[data_w*3 +:data_w];
assign c706ibus[temp_w*4 +:temp_w] = v1858obus[temp_w*1 +:temp_w];
assign v1858ibus[data_w*1 +:data_w] = c706obus[data_w*4 +:data_w];
assign c706ibus[temp_w*5 +:temp_w] = v1954obus[temp_w*0 +:temp_w];
assign v1954ibus[data_w*0 +:data_w] = c706obus[data_w*5 +:data_w];
assign c707ibus[temp_w*0 +:temp_w] = v142obus[temp_w*2 +:temp_w];
assign v142ibus[data_w*2 +:data_w] = c707obus[data_w*0 +:data_w];
assign c707ibus[temp_w*1 +:temp_w] = v204obus[temp_w*4 +:temp_w];
assign v204ibus[data_w*4 +:data_w] = c707obus[data_w*1 +:data_w];
assign c707ibus[temp_w*2 +:temp_w] = v613obus[temp_w*2 +:temp_w];
assign v613ibus[data_w*2 +:data_w] = c707obus[data_w*2 +:data_w];
assign c707ibus[temp_w*3 +:temp_w] = v946obus[temp_w*4 +:temp_w];
assign v946ibus[data_w*4 +:data_w] = c707obus[data_w*3 +:data_w];
assign c707ibus[temp_w*4 +:temp_w] = v1859obus[temp_w*1 +:temp_w];
assign v1859ibus[data_w*1 +:data_w] = c707obus[data_w*4 +:data_w];
assign c707ibus[temp_w*5 +:temp_w] = v1955obus[temp_w*0 +:temp_w];
assign v1955ibus[data_w*0 +:data_w] = c707obus[data_w*5 +:data_w];
assign c708ibus[temp_w*0 +:temp_w] = v143obus[temp_w*2 +:temp_w];
assign v143ibus[data_w*2 +:data_w] = c708obus[data_w*0 +:data_w];
assign c708ibus[temp_w*1 +:temp_w] = v205obus[temp_w*4 +:temp_w];
assign v205ibus[data_w*4 +:data_w] = c708obus[data_w*1 +:data_w];
assign c708ibus[temp_w*2 +:temp_w] = v614obus[temp_w*2 +:temp_w];
assign v614ibus[data_w*2 +:data_w] = c708obus[data_w*2 +:data_w];
assign c708ibus[temp_w*3 +:temp_w] = v947obus[temp_w*4 +:temp_w];
assign v947ibus[data_w*4 +:data_w] = c708obus[data_w*3 +:data_w];
assign c708ibus[temp_w*4 +:temp_w] = v1860obus[temp_w*1 +:temp_w];
assign v1860ibus[data_w*1 +:data_w] = c708obus[data_w*4 +:data_w];
assign c708ibus[temp_w*5 +:temp_w] = v1956obus[temp_w*0 +:temp_w];
assign v1956ibus[data_w*0 +:data_w] = c708obus[data_w*5 +:data_w];
assign c709ibus[temp_w*0 +:temp_w] = v144obus[temp_w*2 +:temp_w];
assign v144ibus[data_w*2 +:data_w] = c709obus[data_w*0 +:data_w];
assign c709ibus[temp_w*1 +:temp_w] = v206obus[temp_w*4 +:temp_w];
assign v206ibus[data_w*4 +:data_w] = c709obus[data_w*1 +:data_w];
assign c709ibus[temp_w*2 +:temp_w] = v615obus[temp_w*2 +:temp_w];
assign v615ibus[data_w*2 +:data_w] = c709obus[data_w*2 +:data_w];
assign c709ibus[temp_w*3 +:temp_w] = v948obus[temp_w*4 +:temp_w];
assign v948ibus[data_w*4 +:data_w] = c709obus[data_w*3 +:data_w];
assign c709ibus[temp_w*4 +:temp_w] = v1861obus[temp_w*1 +:temp_w];
assign v1861ibus[data_w*1 +:data_w] = c709obus[data_w*4 +:data_w];
assign c709ibus[temp_w*5 +:temp_w] = v1957obus[temp_w*0 +:temp_w];
assign v1957ibus[data_w*0 +:data_w] = c709obus[data_w*5 +:data_w];
assign c710ibus[temp_w*0 +:temp_w] = v145obus[temp_w*2 +:temp_w];
assign v145ibus[data_w*2 +:data_w] = c710obus[data_w*0 +:data_w];
assign c710ibus[temp_w*1 +:temp_w] = v207obus[temp_w*4 +:temp_w];
assign v207ibus[data_w*4 +:data_w] = c710obus[data_w*1 +:data_w];
assign c710ibus[temp_w*2 +:temp_w] = v616obus[temp_w*2 +:temp_w];
assign v616ibus[data_w*2 +:data_w] = c710obus[data_w*2 +:data_w];
assign c710ibus[temp_w*3 +:temp_w] = v949obus[temp_w*4 +:temp_w];
assign v949ibus[data_w*4 +:data_w] = c710obus[data_w*3 +:data_w];
assign c710ibus[temp_w*4 +:temp_w] = v1862obus[temp_w*1 +:temp_w];
assign v1862ibus[data_w*1 +:data_w] = c710obus[data_w*4 +:data_w];
assign c710ibus[temp_w*5 +:temp_w] = v1958obus[temp_w*0 +:temp_w];
assign v1958ibus[data_w*0 +:data_w] = c710obus[data_w*5 +:data_w];
assign c711ibus[temp_w*0 +:temp_w] = v146obus[temp_w*2 +:temp_w];
assign v146ibus[data_w*2 +:data_w] = c711obus[data_w*0 +:data_w];
assign c711ibus[temp_w*1 +:temp_w] = v208obus[temp_w*4 +:temp_w];
assign v208ibus[data_w*4 +:data_w] = c711obus[data_w*1 +:data_w];
assign c711ibus[temp_w*2 +:temp_w] = v617obus[temp_w*2 +:temp_w];
assign v617ibus[data_w*2 +:data_w] = c711obus[data_w*2 +:data_w];
assign c711ibus[temp_w*3 +:temp_w] = v950obus[temp_w*4 +:temp_w];
assign v950ibus[data_w*4 +:data_w] = c711obus[data_w*3 +:data_w];
assign c711ibus[temp_w*4 +:temp_w] = v1863obus[temp_w*1 +:temp_w];
assign v1863ibus[data_w*1 +:data_w] = c711obus[data_w*4 +:data_w];
assign c711ibus[temp_w*5 +:temp_w] = v1959obus[temp_w*0 +:temp_w];
assign v1959ibus[data_w*0 +:data_w] = c711obus[data_w*5 +:data_w];
assign c712ibus[temp_w*0 +:temp_w] = v147obus[temp_w*2 +:temp_w];
assign v147ibus[data_w*2 +:data_w] = c712obus[data_w*0 +:data_w];
assign c712ibus[temp_w*1 +:temp_w] = v209obus[temp_w*4 +:temp_w];
assign v209ibus[data_w*4 +:data_w] = c712obus[data_w*1 +:data_w];
assign c712ibus[temp_w*2 +:temp_w] = v618obus[temp_w*2 +:temp_w];
assign v618ibus[data_w*2 +:data_w] = c712obus[data_w*2 +:data_w];
assign c712ibus[temp_w*3 +:temp_w] = v951obus[temp_w*4 +:temp_w];
assign v951ibus[data_w*4 +:data_w] = c712obus[data_w*3 +:data_w];
assign c712ibus[temp_w*4 +:temp_w] = v1864obus[temp_w*1 +:temp_w];
assign v1864ibus[data_w*1 +:data_w] = c712obus[data_w*4 +:data_w];
assign c712ibus[temp_w*5 +:temp_w] = v1960obus[temp_w*0 +:temp_w];
assign v1960ibus[data_w*0 +:data_w] = c712obus[data_w*5 +:data_w];
assign c713ibus[temp_w*0 +:temp_w] = v148obus[temp_w*2 +:temp_w];
assign v148ibus[data_w*2 +:data_w] = c713obus[data_w*0 +:data_w];
assign c713ibus[temp_w*1 +:temp_w] = v210obus[temp_w*4 +:temp_w];
assign v210ibus[data_w*4 +:data_w] = c713obus[data_w*1 +:data_w];
assign c713ibus[temp_w*2 +:temp_w] = v619obus[temp_w*2 +:temp_w];
assign v619ibus[data_w*2 +:data_w] = c713obus[data_w*2 +:data_w];
assign c713ibus[temp_w*3 +:temp_w] = v952obus[temp_w*4 +:temp_w];
assign v952ibus[data_w*4 +:data_w] = c713obus[data_w*3 +:data_w];
assign c713ibus[temp_w*4 +:temp_w] = v1865obus[temp_w*1 +:temp_w];
assign v1865ibus[data_w*1 +:data_w] = c713obus[data_w*4 +:data_w];
assign c713ibus[temp_w*5 +:temp_w] = v1961obus[temp_w*0 +:temp_w];
assign v1961ibus[data_w*0 +:data_w] = c713obus[data_w*5 +:data_w];
assign c714ibus[temp_w*0 +:temp_w] = v149obus[temp_w*2 +:temp_w];
assign v149ibus[data_w*2 +:data_w] = c714obus[data_w*0 +:data_w];
assign c714ibus[temp_w*1 +:temp_w] = v211obus[temp_w*4 +:temp_w];
assign v211ibus[data_w*4 +:data_w] = c714obus[data_w*1 +:data_w];
assign c714ibus[temp_w*2 +:temp_w] = v620obus[temp_w*2 +:temp_w];
assign v620ibus[data_w*2 +:data_w] = c714obus[data_w*2 +:data_w];
assign c714ibus[temp_w*3 +:temp_w] = v953obus[temp_w*4 +:temp_w];
assign v953ibus[data_w*4 +:data_w] = c714obus[data_w*3 +:data_w];
assign c714ibus[temp_w*4 +:temp_w] = v1866obus[temp_w*1 +:temp_w];
assign v1866ibus[data_w*1 +:data_w] = c714obus[data_w*4 +:data_w];
assign c714ibus[temp_w*5 +:temp_w] = v1962obus[temp_w*0 +:temp_w];
assign v1962ibus[data_w*0 +:data_w] = c714obus[data_w*5 +:data_w];
assign c715ibus[temp_w*0 +:temp_w] = v150obus[temp_w*2 +:temp_w];
assign v150ibus[data_w*2 +:data_w] = c715obus[data_w*0 +:data_w];
assign c715ibus[temp_w*1 +:temp_w] = v212obus[temp_w*4 +:temp_w];
assign v212ibus[data_w*4 +:data_w] = c715obus[data_w*1 +:data_w];
assign c715ibus[temp_w*2 +:temp_w] = v621obus[temp_w*2 +:temp_w];
assign v621ibus[data_w*2 +:data_w] = c715obus[data_w*2 +:data_w];
assign c715ibus[temp_w*3 +:temp_w] = v954obus[temp_w*4 +:temp_w];
assign v954ibus[data_w*4 +:data_w] = c715obus[data_w*3 +:data_w];
assign c715ibus[temp_w*4 +:temp_w] = v1867obus[temp_w*1 +:temp_w];
assign v1867ibus[data_w*1 +:data_w] = c715obus[data_w*4 +:data_w];
assign c715ibus[temp_w*5 +:temp_w] = v1963obus[temp_w*0 +:temp_w];
assign v1963ibus[data_w*0 +:data_w] = c715obus[data_w*5 +:data_w];
assign c716ibus[temp_w*0 +:temp_w] = v151obus[temp_w*2 +:temp_w];
assign v151ibus[data_w*2 +:data_w] = c716obus[data_w*0 +:data_w];
assign c716ibus[temp_w*1 +:temp_w] = v213obus[temp_w*4 +:temp_w];
assign v213ibus[data_w*4 +:data_w] = c716obus[data_w*1 +:data_w];
assign c716ibus[temp_w*2 +:temp_w] = v622obus[temp_w*2 +:temp_w];
assign v622ibus[data_w*2 +:data_w] = c716obus[data_w*2 +:data_w];
assign c716ibus[temp_w*3 +:temp_w] = v955obus[temp_w*4 +:temp_w];
assign v955ibus[data_w*4 +:data_w] = c716obus[data_w*3 +:data_w];
assign c716ibus[temp_w*4 +:temp_w] = v1868obus[temp_w*1 +:temp_w];
assign v1868ibus[data_w*1 +:data_w] = c716obus[data_w*4 +:data_w];
assign c716ibus[temp_w*5 +:temp_w] = v1964obus[temp_w*0 +:temp_w];
assign v1964ibus[data_w*0 +:data_w] = c716obus[data_w*5 +:data_w];
assign c717ibus[temp_w*0 +:temp_w] = v152obus[temp_w*2 +:temp_w];
assign v152ibus[data_w*2 +:data_w] = c717obus[data_w*0 +:data_w];
assign c717ibus[temp_w*1 +:temp_w] = v214obus[temp_w*4 +:temp_w];
assign v214ibus[data_w*4 +:data_w] = c717obus[data_w*1 +:data_w];
assign c717ibus[temp_w*2 +:temp_w] = v623obus[temp_w*2 +:temp_w];
assign v623ibus[data_w*2 +:data_w] = c717obus[data_w*2 +:data_w];
assign c717ibus[temp_w*3 +:temp_w] = v956obus[temp_w*4 +:temp_w];
assign v956ibus[data_w*4 +:data_w] = c717obus[data_w*3 +:data_w];
assign c717ibus[temp_w*4 +:temp_w] = v1869obus[temp_w*1 +:temp_w];
assign v1869ibus[data_w*1 +:data_w] = c717obus[data_w*4 +:data_w];
assign c717ibus[temp_w*5 +:temp_w] = v1965obus[temp_w*0 +:temp_w];
assign v1965ibus[data_w*0 +:data_w] = c717obus[data_w*5 +:data_w];
assign c718ibus[temp_w*0 +:temp_w] = v153obus[temp_w*2 +:temp_w];
assign v153ibus[data_w*2 +:data_w] = c718obus[data_w*0 +:data_w];
assign c718ibus[temp_w*1 +:temp_w] = v215obus[temp_w*4 +:temp_w];
assign v215ibus[data_w*4 +:data_w] = c718obus[data_w*1 +:data_w];
assign c718ibus[temp_w*2 +:temp_w] = v624obus[temp_w*2 +:temp_w];
assign v624ibus[data_w*2 +:data_w] = c718obus[data_w*2 +:data_w];
assign c718ibus[temp_w*3 +:temp_w] = v957obus[temp_w*4 +:temp_w];
assign v957ibus[data_w*4 +:data_w] = c718obus[data_w*3 +:data_w];
assign c718ibus[temp_w*4 +:temp_w] = v1870obus[temp_w*1 +:temp_w];
assign v1870ibus[data_w*1 +:data_w] = c718obus[data_w*4 +:data_w];
assign c718ibus[temp_w*5 +:temp_w] = v1966obus[temp_w*0 +:temp_w];
assign v1966ibus[data_w*0 +:data_w] = c718obus[data_w*5 +:data_w];
assign c719ibus[temp_w*0 +:temp_w] = v154obus[temp_w*2 +:temp_w];
assign v154ibus[data_w*2 +:data_w] = c719obus[data_w*0 +:data_w];
assign c719ibus[temp_w*1 +:temp_w] = v216obus[temp_w*4 +:temp_w];
assign v216ibus[data_w*4 +:data_w] = c719obus[data_w*1 +:data_w];
assign c719ibus[temp_w*2 +:temp_w] = v625obus[temp_w*2 +:temp_w];
assign v625ibus[data_w*2 +:data_w] = c719obus[data_w*2 +:data_w];
assign c719ibus[temp_w*3 +:temp_w] = v958obus[temp_w*4 +:temp_w];
assign v958ibus[data_w*4 +:data_w] = c719obus[data_w*3 +:data_w];
assign c719ibus[temp_w*4 +:temp_w] = v1871obus[temp_w*1 +:temp_w];
assign v1871ibus[data_w*1 +:data_w] = c719obus[data_w*4 +:data_w];
assign c719ibus[temp_w*5 +:temp_w] = v1967obus[temp_w*0 +:temp_w];
assign v1967ibus[data_w*0 +:data_w] = c719obus[data_w*5 +:data_w];
assign c720ibus[temp_w*0 +:temp_w] = v155obus[temp_w*2 +:temp_w];
assign v155ibus[data_w*2 +:data_w] = c720obus[data_w*0 +:data_w];
assign c720ibus[temp_w*1 +:temp_w] = v217obus[temp_w*4 +:temp_w];
assign v217ibus[data_w*4 +:data_w] = c720obus[data_w*1 +:data_w];
assign c720ibus[temp_w*2 +:temp_w] = v626obus[temp_w*2 +:temp_w];
assign v626ibus[data_w*2 +:data_w] = c720obus[data_w*2 +:data_w];
assign c720ibus[temp_w*3 +:temp_w] = v959obus[temp_w*4 +:temp_w];
assign v959ibus[data_w*4 +:data_w] = c720obus[data_w*3 +:data_w];
assign c720ibus[temp_w*4 +:temp_w] = v1872obus[temp_w*1 +:temp_w];
assign v1872ibus[data_w*1 +:data_w] = c720obus[data_w*4 +:data_w];
assign c720ibus[temp_w*5 +:temp_w] = v1968obus[temp_w*0 +:temp_w];
assign v1968ibus[data_w*0 +:data_w] = c720obus[data_w*5 +:data_w];
assign c721ibus[temp_w*0 +:temp_w] = v156obus[temp_w*2 +:temp_w];
assign v156ibus[data_w*2 +:data_w] = c721obus[data_w*0 +:data_w];
assign c721ibus[temp_w*1 +:temp_w] = v218obus[temp_w*4 +:temp_w];
assign v218ibus[data_w*4 +:data_w] = c721obus[data_w*1 +:data_w];
assign c721ibus[temp_w*2 +:temp_w] = v627obus[temp_w*2 +:temp_w];
assign v627ibus[data_w*2 +:data_w] = c721obus[data_w*2 +:data_w];
assign c721ibus[temp_w*3 +:temp_w] = v864obus[temp_w*4 +:temp_w];
assign v864ibus[data_w*4 +:data_w] = c721obus[data_w*3 +:data_w];
assign c721ibus[temp_w*4 +:temp_w] = v1873obus[temp_w*1 +:temp_w];
assign v1873ibus[data_w*1 +:data_w] = c721obus[data_w*4 +:data_w];
assign c721ibus[temp_w*5 +:temp_w] = v1969obus[temp_w*0 +:temp_w];
assign v1969ibus[data_w*0 +:data_w] = c721obus[data_w*5 +:data_w];
assign c722ibus[temp_w*0 +:temp_w] = v157obus[temp_w*2 +:temp_w];
assign v157ibus[data_w*2 +:data_w] = c722obus[data_w*0 +:data_w];
assign c722ibus[temp_w*1 +:temp_w] = v219obus[temp_w*4 +:temp_w];
assign v219ibus[data_w*4 +:data_w] = c722obus[data_w*1 +:data_w];
assign c722ibus[temp_w*2 +:temp_w] = v628obus[temp_w*2 +:temp_w];
assign v628ibus[data_w*2 +:data_w] = c722obus[data_w*2 +:data_w];
assign c722ibus[temp_w*3 +:temp_w] = v865obus[temp_w*4 +:temp_w];
assign v865ibus[data_w*4 +:data_w] = c722obus[data_w*3 +:data_w];
assign c722ibus[temp_w*4 +:temp_w] = v1874obus[temp_w*1 +:temp_w];
assign v1874ibus[data_w*1 +:data_w] = c722obus[data_w*4 +:data_w];
assign c722ibus[temp_w*5 +:temp_w] = v1970obus[temp_w*0 +:temp_w];
assign v1970ibus[data_w*0 +:data_w] = c722obus[data_w*5 +:data_w];
assign c723ibus[temp_w*0 +:temp_w] = v158obus[temp_w*2 +:temp_w];
assign v158ibus[data_w*2 +:data_w] = c723obus[data_w*0 +:data_w];
assign c723ibus[temp_w*1 +:temp_w] = v220obus[temp_w*4 +:temp_w];
assign v220ibus[data_w*4 +:data_w] = c723obus[data_w*1 +:data_w];
assign c723ibus[temp_w*2 +:temp_w] = v629obus[temp_w*2 +:temp_w];
assign v629ibus[data_w*2 +:data_w] = c723obus[data_w*2 +:data_w];
assign c723ibus[temp_w*3 +:temp_w] = v866obus[temp_w*4 +:temp_w];
assign v866ibus[data_w*4 +:data_w] = c723obus[data_w*3 +:data_w];
assign c723ibus[temp_w*4 +:temp_w] = v1875obus[temp_w*1 +:temp_w];
assign v1875ibus[data_w*1 +:data_w] = c723obus[data_w*4 +:data_w];
assign c723ibus[temp_w*5 +:temp_w] = v1971obus[temp_w*0 +:temp_w];
assign v1971ibus[data_w*0 +:data_w] = c723obus[data_w*5 +:data_w];
assign c724ibus[temp_w*0 +:temp_w] = v159obus[temp_w*2 +:temp_w];
assign v159ibus[data_w*2 +:data_w] = c724obus[data_w*0 +:data_w];
assign c724ibus[temp_w*1 +:temp_w] = v221obus[temp_w*4 +:temp_w];
assign v221ibus[data_w*4 +:data_w] = c724obus[data_w*1 +:data_w];
assign c724ibus[temp_w*2 +:temp_w] = v630obus[temp_w*2 +:temp_w];
assign v630ibus[data_w*2 +:data_w] = c724obus[data_w*2 +:data_w];
assign c724ibus[temp_w*3 +:temp_w] = v867obus[temp_w*4 +:temp_w];
assign v867ibus[data_w*4 +:data_w] = c724obus[data_w*3 +:data_w];
assign c724ibus[temp_w*4 +:temp_w] = v1876obus[temp_w*1 +:temp_w];
assign v1876ibus[data_w*1 +:data_w] = c724obus[data_w*4 +:data_w];
assign c724ibus[temp_w*5 +:temp_w] = v1972obus[temp_w*0 +:temp_w];
assign v1972ibus[data_w*0 +:data_w] = c724obus[data_w*5 +:data_w];
assign c725ibus[temp_w*0 +:temp_w] = v160obus[temp_w*2 +:temp_w];
assign v160ibus[data_w*2 +:data_w] = c725obus[data_w*0 +:data_w];
assign c725ibus[temp_w*1 +:temp_w] = v222obus[temp_w*4 +:temp_w];
assign v222ibus[data_w*4 +:data_w] = c725obus[data_w*1 +:data_w];
assign c725ibus[temp_w*2 +:temp_w] = v631obus[temp_w*2 +:temp_w];
assign v631ibus[data_w*2 +:data_w] = c725obus[data_w*2 +:data_w];
assign c725ibus[temp_w*3 +:temp_w] = v868obus[temp_w*4 +:temp_w];
assign v868ibus[data_w*4 +:data_w] = c725obus[data_w*3 +:data_w];
assign c725ibus[temp_w*4 +:temp_w] = v1877obus[temp_w*1 +:temp_w];
assign v1877ibus[data_w*1 +:data_w] = c725obus[data_w*4 +:data_w];
assign c725ibus[temp_w*5 +:temp_w] = v1973obus[temp_w*0 +:temp_w];
assign v1973ibus[data_w*0 +:data_w] = c725obus[data_w*5 +:data_w];
assign c726ibus[temp_w*0 +:temp_w] = v161obus[temp_w*2 +:temp_w];
assign v161ibus[data_w*2 +:data_w] = c726obus[data_w*0 +:data_w];
assign c726ibus[temp_w*1 +:temp_w] = v223obus[temp_w*4 +:temp_w];
assign v223ibus[data_w*4 +:data_w] = c726obus[data_w*1 +:data_w];
assign c726ibus[temp_w*2 +:temp_w] = v632obus[temp_w*2 +:temp_w];
assign v632ibus[data_w*2 +:data_w] = c726obus[data_w*2 +:data_w];
assign c726ibus[temp_w*3 +:temp_w] = v869obus[temp_w*4 +:temp_w];
assign v869ibus[data_w*4 +:data_w] = c726obus[data_w*3 +:data_w];
assign c726ibus[temp_w*4 +:temp_w] = v1878obus[temp_w*1 +:temp_w];
assign v1878ibus[data_w*1 +:data_w] = c726obus[data_w*4 +:data_w];
assign c726ibus[temp_w*5 +:temp_w] = v1974obus[temp_w*0 +:temp_w];
assign v1974ibus[data_w*0 +:data_w] = c726obus[data_w*5 +:data_w];
assign c727ibus[temp_w*0 +:temp_w] = v162obus[temp_w*2 +:temp_w];
assign v162ibus[data_w*2 +:data_w] = c727obus[data_w*0 +:data_w];
assign c727ibus[temp_w*1 +:temp_w] = v224obus[temp_w*4 +:temp_w];
assign v224ibus[data_w*4 +:data_w] = c727obus[data_w*1 +:data_w];
assign c727ibus[temp_w*2 +:temp_w] = v633obus[temp_w*2 +:temp_w];
assign v633ibus[data_w*2 +:data_w] = c727obus[data_w*2 +:data_w];
assign c727ibus[temp_w*3 +:temp_w] = v870obus[temp_w*4 +:temp_w];
assign v870ibus[data_w*4 +:data_w] = c727obus[data_w*3 +:data_w];
assign c727ibus[temp_w*4 +:temp_w] = v1879obus[temp_w*1 +:temp_w];
assign v1879ibus[data_w*1 +:data_w] = c727obus[data_w*4 +:data_w];
assign c727ibus[temp_w*5 +:temp_w] = v1975obus[temp_w*0 +:temp_w];
assign v1975ibus[data_w*0 +:data_w] = c727obus[data_w*5 +:data_w];
assign c728ibus[temp_w*0 +:temp_w] = v163obus[temp_w*2 +:temp_w];
assign v163ibus[data_w*2 +:data_w] = c728obus[data_w*0 +:data_w];
assign c728ibus[temp_w*1 +:temp_w] = v225obus[temp_w*4 +:temp_w];
assign v225ibus[data_w*4 +:data_w] = c728obus[data_w*1 +:data_w];
assign c728ibus[temp_w*2 +:temp_w] = v634obus[temp_w*2 +:temp_w];
assign v634ibus[data_w*2 +:data_w] = c728obus[data_w*2 +:data_w];
assign c728ibus[temp_w*3 +:temp_w] = v871obus[temp_w*4 +:temp_w];
assign v871ibus[data_w*4 +:data_w] = c728obus[data_w*3 +:data_w];
assign c728ibus[temp_w*4 +:temp_w] = v1880obus[temp_w*1 +:temp_w];
assign v1880ibus[data_w*1 +:data_w] = c728obus[data_w*4 +:data_w];
assign c728ibus[temp_w*5 +:temp_w] = v1976obus[temp_w*0 +:temp_w];
assign v1976ibus[data_w*0 +:data_w] = c728obus[data_w*5 +:data_w];
assign c729ibus[temp_w*0 +:temp_w] = v164obus[temp_w*2 +:temp_w];
assign v164ibus[data_w*2 +:data_w] = c729obus[data_w*0 +:data_w];
assign c729ibus[temp_w*1 +:temp_w] = v226obus[temp_w*4 +:temp_w];
assign v226ibus[data_w*4 +:data_w] = c729obus[data_w*1 +:data_w];
assign c729ibus[temp_w*2 +:temp_w] = v635obus[temp_w*2 +:temp_w];
assign v635ibus[data_w*2 +:data_w] = c729obus[data_w*2 +:data_w];
assign c729ibus[temp_w*3 +:temp_w] = v872obus[temp_w*4 +:temp_w];
assign v872ibus[data_w*4 +:data_w] = c729obus[data_w*3 +:data_w];
assign c729ibus[temp_w*4 +:temp_w] = v1881obus[temp_w*1 +:temp_w];
assign v1881ibus[data_w*1 +:data_w] = c729obus[data_w*4 +:data_w];
assign c729ibus[temp_w*5 +:temp_w] = v1977obus[temp_w*0 +:temp_w];
assign v1977ibus[data_w*0 +:data_w] = c729obus[data_w*5 +:data_w];
assign c730ibus[temp_w*0 +:temp_w] = v165obus[temp_w*2 +:temp_w];
assign v165ibus[data_w*2 +:data_w] = c730obus[data_w*0 +:data_w];
assign c730ibus[temp_w*1 +:temp_w] = v227obus[temp_w*4 +:temp_w];
assign v227ibus[data_w*4 +:data_w] = c730obus[data_w*1 +:data_w];
assign c730ibus[temp_w*2 +:temp_w] = v636obus[temp_w*2 +:temp_w];
assign v636ibus[data_w*2 +:data_w] = c730obus[data_w*2 +:data_w];
assign c730ibus[temp_w*3 +:temp_w] = v873obus[temp_w*4 +:temp_w];
assign v873ibus[data_w*4 +:data_w] = c730obus[data_w*3 +:data_w];
assign c730ibus[temp_w*4 +:temp_w] = v1882obus[temp_w*1 +:temp_w];
assign v1882ibus[data_w*1 +:data_w] = c730obus[data_w*4 +:data_w];
assign c730ibus[temp_w*5 +:temp_w] = v1978obus[temp_w*0 +:temp_w];
assign v1978ibus[data_w*0 +:data_w] = c730obus[data_w*5 +:data_w];
assign c731ibus[temp_w*0 +:temp_w] = v166obus[temp_w*2 +:temp_w];
assign v166ibus[data_w*2 +:data_w] = c731obus[data_w*0 +:data_w];
assign c731ibus[temp_w*1 +:temp_w] = v228obus[temp_w*4 +:temp_w];
assign v228ibus[data_w*4 +:data_w] = c731obus[data_w*1 +:data_w];
assign c731ibus[temp_w*2 +:temp_w] = v637obus[temp_w*2 +:temp_w];
assign v637ibus[data_w*2 +:data_w] = c731obus[data_w*2 +:data_w];
assign c731ibus[temp_w*3 +:temp_w] = v874obus[temp_w*4 +:temp_w];
assign v874ibus[data_w*4 +:data_w] = c731obus[data_w*3 +:data_w];
assign c731ibus[temp_w*4 +:temp_w] = v1883obus[temp_w*1 +:temp_w];
assign v1883ibus[data_w*1 +:data_w] = c731obus[data_w*4 +:data_w];
assign c731ibus[temp_w*5 +:temp_w] = v1979obus[temp_w*0 +:temp_w];
assign v1979ibus[data_w*0 +:data_w] = c731obus[data_w*5 +:data_w];
assign c732ibus[temp_w*0 +:temp_w] = v167obus[temp_w*2 +:temp_w];
assign v167ibus[data_w*2 +:data_w] = c732obus[data_w*0 +:data_w];
assign c732ibus[temp_w*1 +:temp_w] = v229obus[temp_w*4 +:temp_w];
assign v229ibus[data_w*4 +:data_w] = c732obus[data_w*1 +:data_w];
assign c732ibus[temp_w*2 +:temp_w] = v638obus[temp_w*2 +:temp_w];
assign v638ibus[data_w*2 +:data_w] = c732obus[data_w*2 +:data_w];
assign c732ibus[temp_w*3 +:temp_w] = v875obus[temp_w*4 +:temp_w];
assign v875ibus[data_w*4 +:data_w] = c732obus[data_w*3 +:data_w];
assign c732ibus[temp_w*4 +:temp_w] = v1884obus[temp_w*1 +:temp_w];
assign v1884ibus[data_w*1 +:data_w] = c732obus[data_w*4 +:data_w];
assign c732ibus[temp_w*5 +:temp_w] = v1980obus[temp_w*0 +:temp_w];
assign v1980ibus[data_w*0 +:data_w] = c732obus[data_w*5 +:data_w];
assign c733ibus[temp_w*0 +:temp_w] = v168obus[temp_w*2 +:temp_w];
assign v168ibus[data_w*2 +:data_w] = c733obus[data_w*0 +:data_w];
assign c733ibus[temp_w*1 +:temp_w] = v230obus[temp_w*4 +:temp_w];
assign v230ibus[data_w*4 +:data_w] = c733obus[data_w*1 +:data_w];
assign c733ibus[temp_w*2 +:temp_w] = v639obus[temp_w*2 +:temp_w];
assign v639ibus[data_w*2 +:data_w] = c733obus[data_w*2 +:data_w];
assign c733ibus[temp_w*3 +:temp_w] = v876obus[temp_w*4 +:temp_w];
assign v876ibus[data_w*4 +:data_w] = c733obus[data_w*3 +:data_w];
assign c733ibus[temp_w*4 +:temp_w] = v1885obus[temp_w*1 +:temp_w];
assign v1885ibus[data_w*1 +:data_w] = c733obus[data_w*4 +:data_w];
assign c733ibus[temp_w*5 +:temp_w] = v1981obus[temp_w*0 +:temp_w];
assign v1981ibus[data_w*0 +:data_w] = c733obus[data_w*5 +:data_w];
assign c734ibus[temp_w*0 +:temp_w] = v169obus[temp_w*2 +:temp_w];
assign v169ibus[data_w*2 +:data_w] = c734obus[data_w*0 +:data_w];
assign c734ibus[temp_w*1 +:temp_w] = v231obus[temp_w*4 +:temp_w];
assign v231ibus[data_w*4 +:data_w] = c734obus[data_w*1 +:data_w];
assign c734ibus[temp_w*2 +:temp_w] = v640obus[temp_w*2 +:temp_w];
assign v640ibus[data_w*2 +:data_w] = c734obus[data_w*2 +:data_w];
assign c734ibus[temp_w*3 +:temp_w] = v877obus[temp_w*4 +:temp_w];
assign v877ibus[data_w*4 +:data_w] = c734obus[data_w*3 +:data_w];
assign c734ibus[temp_w*4 +:temp_w] = v1886obus[temp_w*1 +:temp_w];
assign v1886ibus[data_w*1 +:data_w] = c734obus[data_w*4 +:data_w];
assign c734ibus[temp_w*5 +:temp_w] = v1982obus[temp_w*0 +:temp_w];
assign v1982ibus[data_w*0 +:data_w] = c734obus[data_w*5 +:data_w];
assign c735ibus[temp_w*0 +:temp_w] = v170obus[temp_w*2 +:temp_w];
assign v170ibus[data_w*2 +:data_w] = c735obus[data_w*0 +:data_w];
assign c735ibus[temp_w*1 +:temp_w] = v232obus[temp_w*4 +:temp_w];
assign v232ibus[data_w*4 +:data_w] = c735obus[data_w*1 +:data_w];
assign c735ibus[temp_w*2 +:temp_w] = v641obus[temp_w*2 +:temp_w];
assign v641ibus[data_w*2 +:data_w] = c735obus[data_w*2 +:data_w];
assign c735ibus[temp_w*3 +:temp_w] = v878obus[temp_w*4 +:temp_w];
assign v878ibus[data_w*4 +:data_w] = c735obus[data_w*3 +:data_w];
assign c735ibus[temp_w*4 +:temp_w] = v1887obus[temp_w*1 +:temp_w];
assign v1887ibus[data_w*1 +:data_w] = c735obus[data_w*4 +:data_w];
assign c735ibus[temp_w*5 +:temp_w] = v1983obus[temp_w*0 +:temp_w];
assign v1983ibus[data_w*0 +:data_w] = c735obus[data_w*5 +:data_w];
assign c736ibus[temp_w*0 +:temp_w] = v171obus[temp_w*2 +:temp_w];
assign v171ibus[data_w*2 +:data_w] = c736obus[data_w*0 +:data_w];
assign c736ibus[temp_w*1 +:temp_w] = v233obus[temp_w*4 +:temp_w];
assign v233ibus[data_w*4 +:data_w] = c736obus[data_w*1 +:data_w];
assign c736ibus[temp_w*2 +:temp_w] = v642obus[temp_w*2 +:temp_w];
assign v642ibus[data_w*2 +:data_w] = c736obus[data_w*2 +:data_w];
assign c736ibus[temp_w*3 +:temp_w] = v879obus[temp_w*4 +:temp_w];
assign v879ibus[data_w*4 +:data_w] = c736obus[data_w*3 +:data_w];
assign c736ibus[temp_w*4 +:temp_w] = v1888obus[temp_w*1 +:temp_w];
assign v1888ibus[data_w*1 +:data_w] = c736obus[data_w*4 +:data_w];
assign c736ibus[temp_w*5 +:temp_w] = v1984obus[temp_w*0 +:temp_w];
assign v1984ibus[data_w*0 +:data_w] = c736obus[data_w*5 +:data_w];
assign c737ibus[temp_w*0 +:temp_w] = v172obus[temp_w*2 +:temp_w];
assign v172ibus[data_w*2 +:data_w] = c737obus[data_w*0 +:data_w];
assign c737ibus[temp_w*1 +:temp_w] = v234obus[temp_w*4 +:temp_w];
assign v234ibus[data_w*4 +:data_w] = c737obus[data_w*1 +:data_w];
assign c737ibus[temp_w*2 +:temp_w] = v643obus[temp_w*2 +:temp_w];
assign v643ibus[data_w*2 +:data_w] = c737obus[data_w*2 +:data_w];
assign c737ibus[temp_w*3 +:temp_w] = v880obus[temp_w*4 +:temp_w];
assign v880ibus[data_w*4 +:data_w] = c737obus[data_w*3 +:data_w];
assign c737ibus[temp_w*4 +:temp_w] = v1889obus[temp_w*1 +:temp_w];
assign v1889ibus[data_w*1 +:data_w] = c737obus[data_w*4 +:data_w];
assign c737ibus[temp_w*5 +:temp_w] = v1985obus[temp_w*0 +:temp_w];
assign v1985ibus[data_w*0 +:data_w] = c737obus[data_w*5 +:data_w];
assign c738ibus[temp_w*0 +:temp_w] = v173obus[temp_w*2 +:temp_w];
assign v173ibus[data_w*2 +:data_w] = c738obus[data_w*0 +:data_w];
assign c738ibus[temp_w*1 +:temp_w] = v235obus[temp_w*4 +:temp_w];
assign v235ibus[data_w*4 +:data_w] = c738obus[data_w*1 +:data_w];
assign c738ibus[temp_w*2 +:temp_w] = v644obus[temp_w*2 +:temp_w];
assign v644ibus[data_w*2 +:data_w] = c738obus[data_w*2 +:data_w];
assign c738ibus[temp_w*3 +:temp_w] = v881obus[temp_w*4 +:temp_w];
assign v881ibus[data_w*4 +:data_w] = c738obus[data_w*3 +:data_w];
assign c738ibus[temp_w*4 +:temp_w] = v1890obus[temp_w*1 +:temp_w];
assign v1890ibus[data_w*1 +:data_w] = c738obus[data_w*4 +:data_w];
assign c738ibus[temp_w*5 +:temp_w] = v1986obus[temp_w*0 +:temp_w];
assign v1986ibus[data_w*0 +:data_w] = c738obus[data_w*5 +:data_w];
assign c739ibus[temp_w*0 +:temp_w] = v174obus[temp_w*2 +:temp_w];
assign v174ibus[data_w*2 +:data_w] = c739obus[data_w*0 +:data_w];
assign c739ibus[temp_w*1 +:temp_w] = v236obus[temp_w*4 +:temp_w];
assign v236ibus[data_w*4 +:data_w] = c739obus[data_w*1 +:data_w];
assign c739ibus[temp_w*2 +:temp_w] = v645obus[temp_w*2 +:temp_w];
assign v645ibus[data_w*2 +:data_w] = c739obus[data_w*2 +:data_w];
assign c739ibus[temp_w*3 +:temp_w] = v882obus[temp_w*4 +:temp_w];
assign v882ibus[data_w*4 +:data_w] = c739obus[data_w*3 +:data_w];
assign c739ibus[temp_w*4 +:temp_w] = v1891obus[temp_w*1 +:temp_w];
assign v1891ibus[data_w*1 +:data_w] = c739obus[data_w*4 +:data_w];
assign c739ibus[temp_w*5 +:temp_w] = v1987obus[temp_w*0 +:temp_w];
assign v1987ibus[data_w*0 +:data_w] = c739obus[data_w*5 +:data_w];
assign c740ibus[temp_w*0 +:temp_w] = v175obus[temp_w*2 +:temp_w];
assign v175ibus[data_w*2 +:data_w] = c740obus[data_w*0 +:data_w];
assign c740ibus[temp_w*1 +:temp_w] = v237obus[temp_w*4 +:temp_w];
assign v237ibus[data_w*4 +:data_w] = c740obus[data_w*1 +:data_w];
assign c740ibus[temp_w*2 +:temp_w] = v646obus[temp_w*2 +:temp_w];
assign v646ibus[data_w*2 +:data_w] = c740obus[data_w*2 +:data_w];
assign c740ibus[temp_w*3 +:temp_w] = v883obus[temp_w*4 +:temp_w];
assign v883ibus[data_w*4 +:data_w] = c740obus[data_w*3 +:data_w];
assign c740ibus[temp_w*4 +:temp_w] = v1892obus[temp_w*1 +:temp_w];
assign v1892ibus[data_w*1 +:data_w] = c740obus[data_w*4 +:data_w];
assign c740ibus[temp_w*5 +:temp_w] = v1988obus[temp_w*0 +:temp_w];
assign v1988ibus[data_w*0 +:data_w] = c740obus[data_w*5 +:data_w];
assign c741ibus[temp_w*0 +:temp_w] = v176obus[temp_w*2 +:temp_w];
assign v176ibus[data_w*2 +:data_w] = c741obus[data_w*0 +:data_w];
assign c741ibus[temp_w*1 +:temp_w] = v238obus[temp_w*4 +:temp_w];
assign v238ibus[data_w*4 +:data_w] = c741obus[data_w*1 +:data_w];
assign c741ibus[temp_w*2 +:temp_w] = v647obus[temp_w*2 +:temp_w];
assign v647ibus[data_w*2 +:data_w] = c741obus[data_w*2 +:data_w];
assign c741ibus[temp_w*3 +:temp_w] = v884obus[temp_w*4 +:temp_w];
assign v884ibus[data_w*4 +:data_w] = c741obus[data_w*3 +:data_w];
assign c741ibus[temp_w*4 +:temp_w] = v1893obus[temp_w*1 +:temp_w];
assign v1893ibus[data_w*1 +:data_w] = c741obus[data_w*4 +:data_w];
assign c741ibus[temp_w*5 +:temp_w] = v1989obus[temp_w*0 +:temp_w];
assign v1989ibus[data_w*0 +:data_w] = c741obus[data_w*5 +:data_w];
assign c742ibus[temp_w*0 +:temp_w] = v177obus[temp_w*2 +:temp_w];
assign v177ibus[data_w*2 +:data_w] = c742obus[data_w*0 +:data_w];
assign c742ibus[temp_w*1 +:temp_w] = v239obus[temp_w*4 +:temp_w];
assign v239ibus[data_w*4 +:data_w] = c742obus[data_w*1 +:data_w];
assign c742ibus[temp_w*2 +:temp_w] = v648obus[temp_w*2 +:temp_w];
assign v648ibus[data_w*2 +:data_w] = c742obus[data_w*2 +:data_w];
assign c742ibus[temp_w*3 +:temp_w] = v885obus[temp_w*4 +:temp_w];
assign v885ibus[data_w*4 +:data_w] = c742obus[data_w*3 +:data_w];
assign c742ibus[temp_w*4 +:temp_w] = v1894obus[temp_w*1 +:temp_w];
assign v1894ibus[data_w*1 +:data_w] = c742obus[data_w*4 +:data_w];
assign c742ibus[temp_w*5 +:temp_w] = v1990obus[temp_w*0 +:temp_w];
assign v1990ibus[data_w*0 +:data_w] = c742obus[data_w*5 +:data_w];
assign c743ibus[temp_w*0 +:temp_w] = v178obus[temp_w*2 +:temp_w];
assign v178ibus[data_w*2 +:data_w] = c743obus[data_w*0 +:data_w];
assign c743ibus[temp_w*1 +:temp_w] = v240obus[temp_w*4 +:temp_w];
assign v240ibus[data_w*4 +:data_w] = c743obus[data_w*1 +:data_w];
assign c743ibus[temp_w*2 +:temp_w] = v649obus[temp_w*2 +:temp_w];
assign v649ibus[data_w*2 +:data_w] = c743obus[data_w*2 +:data_w];
assign c743ibus[temp_w*3 +:temp_w] = v886obus[temp_w*4 +:temp_w];
assign v886ibus[data_w*4 +:data_w] = c743obus[data_w*3 +:data_w];
assign c743ibus[temp_w*4 +:temp_w] = v1895obus[temp_w*1 +:temp_w];
assign v1895ibus[data_w*1 +:data_w] = c743obus[data_w*4 +:data_w];
assign c743ibus[temp_w*5 +:temp_w] = v1991obus[temp_w*0 +:temp_w];
assign v1991ibus[data_w*0 +:data_w] = c743obus[data_w*5 +:data_w];
assign c744ibus[temp_w*0 +:temp_w] = v179obus[temp_w*2 +:temp_w];
assign v179ibus[data_w*2 +:data_w] = c744obus[data_w*0 +:data_w];
assign c744ibus[temp_w*1 +:temp_w] = v241obus[temp_w*4 +:temp_w];
assign v241ibus[data_w*4 +:data_w] = c744obus[data_w*1 +:data_w];
assign c744ibus[temp_w*2 +:temp_w] = v650obus[temp_w*2 +:temp_w];
assign v650ibus[data_w*2 +:data_w] = c744obus[data_w*2 +:data_w];
assign c744ibus[temp_w*3 +:temp_w] = v887obus[temp_w*4 +:temp_w];
assign v887ibus[data_w*4 +:data_w] = c744obus[data_w*3 +:data_w];
assign c744ibus[temp_w*4 +:temp_w] = v1896obus[temp_w*1 +:temp_w];
assign v1896ibus[data_w*1 +:data_w] = c744obus[data_w*4 +:data_w];
assign c744ibus[temp_w*5 +:temp_w] = v1992obus[temp_w*0 +:temp_w];
assign v1992ibus[data_w*0 +:data_w] = c744obus[data_w*5 +:data_w];
assign c745ibus[temp_w*0 +:temp_w] = v180obus[temp_w*2 +:temp_w];
assign v180ibus[data_w*2 +:data_w] = c745obus[data_w*0 +:data_w];
assign c745ibus[temp_w*1 +:temp_w] = v242obus[temp_w*4 +:temp_w];
assign v242ibus[data_w*4 +:data_w] = c745obus[data_w*1 +:data_w];
assign c745ibus[temp_w*2 +:temp_w] = v651obus[temp_w*2 +:temp_w];
assign v651ibus[data_w*2 +:data_w] = c745obus[data_w*2 +:data_w];
assign c745ibus[temp_w*3 +:temp_w] = v888obus[temp_w*4 +:temp_w];
assign v888ibus[data_w*4 +:data_w] = c745obus[data_w*3 +:data_w];
assign c745ibus[temp_w*4 +:temp_w] = v1897obus[temp_w*1 +:temp_w];
assign v1897ibus[data_w*1 +:data_w] = c745obus[data_w*4 +:data_w];
assign c745ibus[temp_w*5 +:temp_w] = v1993obus[temp_w*0 +:temp_w];
assign v1993ibus[data_w*0 +:data_w] = c745obus[data_w*5 +:data_w];
assign c746ibus[temp_w*0 +:temp_w] = v181obus[temp_w*2 +:temp_w];
assign v181ibus[data_w*2 +:data_w] = c746obus[data_w*0 +:data_w];
assign c746ibus[temp_w*1 +:temp_w] = v243obus[temp_w*4 +:temp_w];
assign v243ibus[data_w*4 +:data_w] = c746obus[data_w*1 +:data_w];
assign c746ibus[temp_w*2 +:temp_w] = v652obus[temp_w*2 +:temp_w];
assign v652ibus[data_w*2 +:data_w] = c746obus[data_w*2 +:data_w];
assign c746ibus[temp_w*3 +:temp_w] = v889obus[temp_w*4 +:temp_w];
assign v889ibus[data_w*4 +:data_w] = c746obus[data_w*3 +:data_w];
assign c746ibus[temp_w*4 +:temp_w] = v1898obus[temp_w*1 +:temp_w];
assign v1898ibus[data_w*1 +:data_w] = c746obus[data_w*4 +:data_w];
assign c746ibus[temp_w*5 +:temp_w] = v1994obus[temp_w*0 +:temp_w];
assign v1994ibus[data_w*0 +:data_w] = c746obus[data_w*5 +:data_w];
assign c747ibus[temp_w*0 +:temp_w] = v182obus[temp_w*2 +:temp_w];
assign v182ibus[data_w*2 +:data_w] = c747obus[data_w*0 +:data_w];
assign c747ibus[temp_w*1 +:temp_w] = v244obus[temp_w*4 +:temp_w];
assign v244ibus[data_w*4 +:data_w] = c747obus[data_w*1 +:data_w];
assign c747ibus[temp_w*2 +:temp_w] = v653obus[temp_w*2 +:temp_w];
assign v653ibus[data_w*2 +:data_w] = c747obus[data_w*2 +:data_w];
assign c747ibus[temp_w*3 +:temp_w] = v890obus[temp_w*4 +:temp_w];
assign v890ibus[data_w*4 +:data_w] = c747obus[data_w*3 +:data_w];
assign c747ibus[temp_w*4 +:temp_w] = v1899obus[temp_w*1 +:temp_w];
assign v1899ibus[data_w*1 +:data_w] = c747obus[data_w*4 +:data_w];
assign c747ibus[temp_w*5 +:temp_w] = v1995obus[temp_w*0 +:temp_w];
assign v1995ibus[data_w*0 +:data_w] = c747obus[data_w*5 +:data_w];
assign c748ibus[temp_w*0 +:temp_w] = v183obus[temp_w*2 +:temp_w];
assign v183ibus[data_w*2 +:data_w] = c748obus[data_w*0 +:data_w];
assign c748ibus[temp_w*1 +:temp_w] = v245obus[temp_w*4 +:temp_w];
assign v245ibus[data_w*4 +:data_w] = c748obus[data_w*1 +:data_w];
assign c748ibus[temp_w*2 +:temp_w] = v654obus[temp_w*2 +:temp_w];
assign v654ibus[data_w*2 +:data_w] = c748obus[data_w*2 +:data_w];
assign c748ibus[temp_w*3 +:temp_w] = v891obus[temp_w*4 +:temp_w];
assign v891ibus[data_w*4 +:data_w] = c748obus[data_w*3 +:data_w];
assign c748ibus[temp_w*4 +:temp_w] = v1900obus[temp_w*1 +:temp_w];
assign v1900ibus[data_w*1 +:data_w] = c748obus[data_w*4 +:data_w];
assign c748ibus[temp_w*5 +:temp_w] = v1996obus[temp_w*0 +:temp_w];
assign v1996ibus[data_w*0 +:data_w] = c748obus[data_w*5 +:data_w];
assign c749ibus[temp_w*0 +:temp_w] = v184obus[temp_w*2 +:temp_w];
assign v184ibus[data_w*2 +:data_w] = c749obus[data_w*0 +:data_w];
assign c749ibus[temp_w*1 +:temp_w] = v246obus[temp_w*4 +:temp_w];
assign v246ibus[data_w*4 +:data_w] = c749obus[data_w*1 +:data_w];
assign c749ibus[temp_w*2 +:temp_w] = v655obus[temp_w*2 +:temp_w];
assign v655ibus[data_w*2 +:data_w] = c749obus[data_w*2 +:data_w];
assign c749ibus[temp_w*3 +:temp_w] = v892obus[temp_w*4 +:temp_w];
assign v892ibus[data_w*4 +:data_w] = c749obus[data_w*3 +:data_w];
assign c749ibus[temp_w*4 +:temp_w] = v1901obus[temp_w*1 +:temp_w];
assign v1901ibus[data_w*1 +:data_w] = c749obus[data_w*4 +:data_w];
assign c749ibus[temp_w*5 +:temp_w] = v1997obus[temp_w*0 +:temp_w];
assign v1997ibus[data_w*0 +:data_w] = c749obus[data_w*5 +:data_w];
assign c750ibus[temp_w*0 +:temp_w] = v185obus[temp_w*2 +:temp_w];
assign v185ibus[data_w*2 +:data_w] = c750obus[data_w*0 +:data_w];
assign c750ibus[temp_w*1 +:temp_w] = v247obus[temp_w*4 +:temp_w];
assign v247ibus[data_w*4 +:data_w] = c750obus[data_w*1 +:data_w];
assign c750ibus[temp_w*2 +:temp_w] = v656obus[temp_w*2 +:temp_w];
assign v656ibus[data_w*2 +:data_w] = c750obus[data_w*2 +:data_w];
assign c750ibus[temp_w*3 +:temp_w] = v893obus[temp_w*4 +:temp_w];
assign v893ibus[data_w*4 +:data_w] = c750obus[data_w*3 +:data_w];
assign c750ibus[temp_w*4 +:temp_w] = v1902obus[temp_w*1 +:temp_w];
assign v1902ibus[data_w*1 +:data_w] = c750obus[data_w*4 +:data_w];
assign c750ibus[temp_w*5 +:temp_w] = v1998obus[temp_w*0 +:temp_w];
assign v1998ibus[data_w*0 +:data_w] = c750obus[data_w*5 +:data_w];
assign c751ibus[temp_w*0 +:temp_w] = v186obus[temp_w*2 +:temp_w];
assign v186ibus[data_w*2 +:data_w] = c751obus[data_w*0 +:data_w];
assign c751ibus[temp_w*1 +:temp_w] = v248obus[temp_w*4 +:temp_w];
assign v248ibus[data_w*4 +:data_w] = c751obus[data_w*1 +:data_w];
assign c751ibus[temp_w*2 +:temp_w] = v657obus[temp_w*2 +:temp_w];
assign v657ibus[data_w*2 +:data_w] = c751obus[data_w*2 +:data_w];
assign c751ibus[temp_w*3 +:temp_w] = v894obus[temp_w*4 +:temp_w];
assign v894ibus[data_w*4 +:data_w] = c751obus[data_w*3 +:data_w];
assign c751ibus[temp_w*4 +:temp_w] = v1903obus[temp_w*1 +:temp_w];
assign v1903ibus[data_w*1 +:data_w] = c751obus[data_w*4 +:data_w];
assign c751ibus[temp_w*5 +:temp_w] = v1999obus[temp_w*0 +:temp_w];
assign v1999ibus[data_w*0 +:data_w] = c751obus[data_w*5 +:data_w];
assign c752ibus[temp_w*0 +:temp_w] = v187obus[temp_w*2 +:temp_w];
assign v187ibus[data_w*2 +:data_w] = c752obus[data_w*0 +:data_w];
assign c752ibus[temp_w*1 +:temp_w] = v249obus[temp_w*4 +:temp_w];
assign v249ibus[data_w*4 +:data_w] = c752obus[data_w*1 +:data_w];
assign c752ibus[temp_w*2 +:temp_w] = v658obus[temp_w*2 +:temp_w];
assign v658ibus[data_w*2 +:data_w] = c752obus[data_w*2 +:data_w];
assign c752ibus[temp_w*3 +:temp_w] = v895obus[temp_w*4 +:temp_w];
assign v895ibus[data_w*4 +:data_w] = c752obus[data_w*3 +:data_w];
assign c752ibus[temp_w*4 +:temp_w] = v1904obus[temp_w*1 +:temp_w];
assign v1904ibus[data_w*1 +:data_w] = c752obus[data_w*4 +:data_w];
assign c752ibus[temp_w*5 +:temp_w] = v2000obus[temp_w*0 +:temp_w];
assign v2000ibus[data_w*0 +:data_w] = c752obus[data_w*5 +:data_w];
assign c753ibus[temp_w*0 +:temp_w] = v188obus[temp_w*2 +:temp_w];
assign v188ibus[data_w*2 +:data_w] = c753obus[data_w*0 +:data_w];
assign c753ibus[temp_w*1 +:temp_w] = v250obus[temp_w*4 +:temp_w];
assign v250ibus[data_w*4 +:data_w] = c753obus[data_w*1 +:data_w];
assign c753ibus[temp_w*2 +:temp_w] = v659obus[temp_w*2 +:temp_w];
assign v659ibus[data_w*2 +:data_w] = c753obus[data_w*2 +:data_w];
assign c753ibus[temp_w*3 +:temp_w] = v896obus[temp_w*4 +:temp_w];
assign v896ibus[data_w*4 +:data_w] = c753obus[data_w*3 +:data_w];
assign c753ibus[temp_w*4 +:temp_w] = v1905obus[temp_w*1 +:temp_w];
assign v1905ibus[data_w*1 +:data_w] = c753obus[data_w*4 +:data_w];
assign c753ibus[temp_w*5 +:temp_w] = v2001obus[temp_w*0 +:temp_w];
assign v2001ibus[data_w*0 +:data_w] = c753obus[data_w*5 +:data_w];
assign c754ibus[temp_w*0 +:temp_w] = v189obus[temp_w*2 +:temp_w];
assign v189ibus[data_w*2 +:data_w] = c754obus[data_w*0 +:data_w];
assign c754ibus[temp_w*1 +:temp_w] = v251obus[temp_w*4 +:temp_w];
assign v251ibus[data_w*4 +:data_w] = c754obus[data_w*1 +:data_w];
assign c754ibus[temp_w*2 +:temp_w] = v660obus[temp_w*2 +:temp_w];
assign v660ibus[data_w*2 +:data_w] = c754obus[data_w*2 +:data_w];
assign c754ibus[temp_w*3 +:temp_w] = v897obus[temp_w*4 +:temp_w];
assign v897ibus[data_w*4 +:data_w] = c754obus[data_w*3 +:data_w];
assign c754ibus[temp_w*4 +:temp_w] = v1906obus[temp_w*1 +:temp_w];
assign v1906ibus[data_w*1 +:data_w] = c754obus[data_w*4 +:data_w];
assign c754ibus[temp_w*5 +:temp_w] = v2002obus[temp_w*0 +:temp_w];
assign v2002ibus[data_w*0 +:data_w] = c754obus[data_w*5 +:data_w];
assign c755ibus[temp_w*0 +:temp_w] = v190obus[temp_w*2 +:temp_w];
assign v190ibus[data_w*2 +:data_w] = c755obus[data_w*0 +:data_w];
assign c755ibus[temp_w*1 +:temp_w] = v252obus[temp_w*4 +:temp_w];
assign v252ibus[data_w*4 +:data_w] = c755obus[data_w*1 +:data_w];
assign c755ibus[temp_w*2 +:temp_w] = v661obus[temp_w*2 +:temp_w];
assign v661ibus[data_w*2 +:data_w] = c755obus[data_w*2 +:data_w];
assign c755ibus[temp_w*3 +:temp_w] = v898obus[temp_w*4 +:temp_w];
assign v898ibus[data_w*4 +:data_w] = c755obus[data_w*3 +:data_w];
assign c755ibus[temp_w*4 +:temp_w] = v1907obus[temp_w*1 +:temp_w];
assign v1907ibus[data_w*1 +:data_w] = c755obus[data_w*4 +:data_w];
assign c755ibus[temp_w*5 +:temp_w] = v2003obus[temp_w*0 +:temp_w];
assign v2003ibus[data_w*0 +:data_w] = c755obus[data_w*5 +:data_w];
assign c756ibus[temp_w*0 +:temp_w] = v191obus[temp_w*2 +:temp_w];
assign v191ibus[data_w*2 +:data_w] = c756obus[data_w*0 +:data_w];
assign c756ibus[temp_w*1 +:temp_w] = v253obus[temp_w*4 +:temp_w];
assign v253ibus[data_w*4 +:data_w] = c756obus[data_w*1 +:data_w];
assign c756ibus[temp_w*2 +:temp_w] = v662obus[temp_w*2 +:temp_w];
assign v662ibus[data_w*2 +:data_w] = c756obus[data_w*2 +:data_w];
assign c756ibus[temp_w*3 +:temp_w] = v899obus[temp_w*4 +:temp_w];
assign v899ibus[data_w*4 +:data_w] = c756obus[data_w*3 +:data_w];
assign c756ibus[temp_w*4 +:temp_w] = v1908obus[temp_w*1 +:temp_w];
assign v1908ibus[data_w*1 +:data_w] = c756obus[data_w*4 +:data_w];
assign c756ibus[temp_w*5 +:temp_w] = v2004obus[temp_w*0 +:temp_w];
assign v2004ibus[data_w*0 +:data_w] = c756obus[data_w*5 +:data_w];
assign c757ibus[temp_w*0 +:temp_w] = v96obus[temp_w*2 +:temp_w];
assign v96ibus[data_w*2 +:data_w] = c757obus[data_w*0 +:data_w];
assign c757ibus[temp_w*1 +:temp_w] = v254obus[temp_w*4 +:temp_w];
assign v254ibus[data_w*4 +:data_w] = c757obus[data_w*1 +:data_w];
assign c757ibus[temp_w*2 +:temp_w] = v663obus[temp_w*2 +:temp_w];
assign v663ibus[data_w*2 +:data_w] = c757obus[data_w*2 +:data_w];
assign c757ibus[temp_w*3 +:temp_w] = v900obus[temp_w*4 +:temp_w];
assign v900ibus[data_w*4 +:data_w] = c757obus[data_w*3 +:data_w];
assign c757ibus[temp_w*4 +:temp_w] = v1909obus[temp_w*1 +:temp_w];
assign v1909ibus[data_w*1 +:data_w] = c757obus[data_w*4 +:data_w];
assign c757ibus[temp_w*5 +:temp_w] = v2005obus[temp_w*0 +:temp_w];
assign v2005ibus[data_w*0 +:data_w] = c757obus[data_w*5 +:data_w];
assign c758ibus[temp_w*0 +:temp_w] = v97obus[temp_w*2 +:temp_w];
assign v97ibus[data_w*2 +:data_w] = c758obus[data_w*0 +:data_w];
assign c758ibus[temp_w*1 +:temp_w] = v255obus[temp_w*4 +:temp_w];
assign v255ibus[data_w*4 +:data_w] = c758obus[data_w*1 +:data_w];
assign c758ibus[temp_w*2 +:temp_w] = v664obus[temp_w*2 +:temp_w];
assign v664ibus[data_w*2 +:data_w] = c758obus[data_w*2 +:data_w];
assign c758ibus[temp_w*3 +:temp_w] = v901obus[temp_w*4 +:temp_w];
assign v901ibus[data_w*4 +:data_w] = c758obus[data_w*3 +:data_w];
assign c758ibus[temp_w*4 +:temp_w] = v1910obus[temp_w*1 +:temp_w];
assign v1910ibus[data_w*1 +:data_w] = c758obus[data_w*4 +:data_w];
assign c758ibus[temp_w*5 +:temp_w] = v2006obus[temp_w*0 +:temp_w];
assign v2006ibus[data_w*0 +:data_w] = c758obus[data_w*5 +:data_w];
assign c759ibus[temp_w*0 +:temp_w] = v98obus[temp_w*2 +:temp_w];
assign v98ibus[data_w*2 +:data_w] = c759obus[data_w*0 +:data_w];
assign c759ibus[temp_w*1 +:temp_w] = v256obus[temp_w*4 +:temp_w];
assign v256ibus[data_w*4 +:data_w] = c759obus[data_w*1 +:data_w];
assign c759ibus[temp_w*2 +:temp_w] = v665obus[temp_w*2 +:temp_w];
assign v665ibus[data_w*2 +:data_w] = c759obus[data_w*2 +:data_w];
assign c759ibus[temp_w*3 +:temp_w] = v902obus[temp_w*4 +:temp_w];
assign v902ibus[data_w*4 +:data_w] = c759obus[data_w*3 +:data_w];
assign c759ibus[temp_w*4 +:temp_w] = v1911obus[temp_w*1 +:temp_w];
assign v1911ibus[data_w*1 +:data_w] = c759obus[data_w*4 +:data_w];
assign c759ibus[temp_w*5 +:temp_w] = v2007obus[temp_w*0 +:temp_w];
assign v2007ibus[data_w*0 +:data_w] = c759obus[data_w*5 +:data_w];
assign c760ibus[temp_w*0 +:temp_w] = v99obus[temp_w*2 +:temp_w];
assign v99ibus[data_w*2 +:data_w] = c760obus[data_w*0 +:data_w];
assign c760ibus[temp_w*1 +:temp_w] = v257obus[temp_w*4 +:temp_w];
assign v257ibus[data_w*4 +:data_w] = c760obus[data_w*1 +:data_w];
assign c760ibus[temp_w*2 +:temp_w] = v666obus[temp_w*2 +:temp_w];
assign v666ibus[data_w*2 +:data_w] = c760obus[data_w*2 +:data_w];
assign c760ibus[temp_w*3 +:temp_w] = v903obus[temp_w*4 +:temp_w];
assign v903ibus[data_w*4 +:data_w] = c760obus[data_w*3 +:data_w];
assign c760ibus[temp_w*4 +:temp_w] = v1912obus[temp_w*1 +:temp_w];
assign v1912ibus[data_w*1 +:data_w] = c760obus[data_w*4 +:data_w];
assign c760ibus[temp_w*5 +:temp_w] = v2008obus[temp_w*0 +:temp_w];
assign v2008ibus[data_w*0 +:data_w] = c760obus[data_w*5 +:data_w];
assign c761ibus[temp_w*0 +:temp_w] = v100obus[temp_w*2 +:temp_w];
assign v100ibus[data_w*2 +:data_w] = c761obus[data_w*0 +:data_w];
assign c761ibus[temp_w*1 +:temp_w] = v258obus[temp_w*4 +:temp_w];
assign v258ibus[data_w*4 +:data_w] = c761obus[data_w*1 +:data_w];
assign c761ibus[temp_w*2 +:temp_w] = v667obus[temp_w*2 +:temp_w];
assign v667ibus[data_w*2 +:data_w] = c761obus[data_w*2 +:data_w];
assign c761ibus[temp_w*3 +:temp_w] = v904obus[temp_w*4 +:temp_w];
assign v904ibus[data_w*4 +:data_w] = c761obus[data_w*3 +:data_w];
assign c761ibus[temp_w*4 +:temp_w] = v1913obus[temp_w*1 +:temp_w];
assign v1913ibus[data_w*1 +:data_w] = c761obus[data_w*4 +:data_w];
assign c761ibus[temp_w*5 +:temp_w] = v2009obus[temp_w*0 +:temp_w];
assign v2009ibus[data_w*0 +:data_w] = c761obus[data_w*5 +:data_w];
assign c762ibus[temp_w*0 +:temp_w] = v101obus[temp_w*2 +:temp_w];
assign v101ibus[data_w*2 +:data_w] = c762obus[data_w*0 +:data_w];
assign c762ibus[temp_w*1 +:temp_w] = v259obus[temp_w*4 +:temp_w];
assign v259ibus[data_w*4 +:data_w] = c762obus[data_w*1 +:data_w];
assign c762ibus[temp_w*2 +:temp_w] = v668obus[temp_w*2 +:temp_w];
assign v668ibus[data_w*2 +:data_w] = c762obus[data_w*2 +:data_w];
assign c762ibus[temp_w*3 +:temp_w] = v905obus[temp_w*4 +:temp_w];
assign v905ibus[data_w*4 +:data_w] = c762obus[data_w*3 +:data_w];
assign c762ibus[temp_w*4 +:temp_w] = v1914obus[temp_w*1 +:temp_w];
assign v1914ibus[data_w*1 +:data_w] = c762obus[data_w*4 +:data_w];
assign c762ibus[temp_w*5 +:temp_w] = v2010obus[temp_w*0 +:temp_w];
assign v2010ibus[data_w*0 +:data_w] = c762obus[data_w*5 +:data_w];
assign c763ibus[temp_w*0 +:temp_w] = v102obus[temp_w*2 +:temp_w];
assign v102ibus[data_w*2 +:data_w] = c763obus[data_w*0 +:data_w];
assign c763ibus[temp_w*1 +:temp_w] = v260obus[temp_w*4 +:temp_w];
assign v260ibus[data_w*4 +:data_w] = c763obus[data_w*1 +:data_w];
assign c763ibus[temp_w*2 +:temp_w] = v669obus[temp_w*2 +:temp_w];
assign v669ibus[data_w*2 +:data_w] = c763obus[data_w*2 +:data_w];
assign c763ibus[temp_w*3 +:temp_w] = v906obus[temp_w*4 +:temp_w];
assign v906ibus[data_w*4 +:data_w] = c763obus[data_w*3 +:data_w];
assign c763ibus[temp_w*4 +:temp_w] = v1915obus[temp_w*1 +:temp_w];
assign v1915ibus[data_w*1 +:data_w] = c763obus[data_w*4 +:data_w];
assign c763ibus[temp_w*5 +:temp_w] = v2011obus[temp_w*0 +:temp_w];
assign v2011ibus[data_w*0 +:data_w] = c763obus[data_w*5 +:data_w];
assign c764ibus[temp_w*0 +:temp_w] = v103obus[temp_w*2 +:temp_w];
assign v103ibus[data_w*2 +:data_w] = c764obus[data_w*0 +:data_w];
assign c764ibus[temp_w*1 +:temp_w] = v261obus[temp_w*4 +:temp_w];
assign v261ibus[data_w*4 +:data_w] = c764obus[data_w*1 +:data_w];
assign c764ibus[temp_w*2 +:temp_w] = v670obus[temp_w*2 +:temp_w];
assign v670ibus[data_w*2 +:data_w] = c764obus[data_w*2 +:data_w];
assign c764ibus[temp_w*3 +:temp_w] = v907obus[temp_w*4 +:temp_w];
assign v907ibus[data_w*4 +:data_w] = c764obus[data_w*3 +:data_w];
assign c764ibus[temp_w*4 +:temp_w] = v1916obus[temp_w*1 +:temp_w];
assign v1916ibus[data_w*1 +:data_w] = c764obus[data_w*4 +:data_w];
assign c764ibus[temp_w*5 +:temp_w] = v2012obus[temp_w*0 +:temp_w];
assign v2012ibus[data_w*0 +:data_w] = c764obus[data_w*5 +:data_w];
assign c765ibus[temp_w*0 +:temp_w] = v104obus[temp_w*2 +:temp_w];
assign v104ibus[data_w*2 +:data_w] = c765obus[data_w*0 +:data_w];
assign c765ibus[temp_w*1 +:temp_w] = v262obus[temp_w*4 +:temp_w];
assign v262ibus[data_w*4 +:data_w] = c765obus[data_w*1 +:data_w];
assign c765ibus[temp_w*2 +:temp_w] = v671obus[temp_w*2 +:temp_w];
assign v671ibus[data_w*2 +:data_w] = c765obus[data_w*2 +:data_w];
assign c765ibus[temp_w*3 +:temp_w] = v908obus[temp_w*4 +:temp_w];
assign v908ibus[data_w*4 +:data_w] = c765obus[data_w*3 +:data_w];
assign c765ibus[temp_w*4 +:temp_w] = v1917obus[temp_w*1 +:temp_w];
assign v1917ibus[data_w*1 +:data_w] = c765obus[data_w*4 +:data_w];
assign c765ibus[temp_w*5 +:temp_w] = v2013obus[temp_w*0 +:temp_w];
assign v2013ibus[data_w*0 +:data_w] = c765obus[data_w*5 +:data_w];
assign c766ibus[temp_w*0 +:temp_w] = v105obus[temp_w*2 +:temp_w];
assign v105ibus[data_w*2 +:data_w] = c766obus[data_w*0 +:data_w];
assign c766ibus[temp_w*1 +:temp_w] = v263obus[temp_w*4 +:temp_w];
assign v263ibus[data_w*4 +:data_w] = c766obus[data_w*1 +:data_w];
assign c766ibus[temp_w*2 +:temp_w] = v576obus[temp_w*2 +:temp_w];
assign v576ibus[data_w*2 +:data_w] = c766obus[data_w*2 +:data_w];
assign c766ibus[temp_w*3 +:temp_w] = v909obus[temp_w*4 +:temp_w];
assign v909ibus[data_w*4 +:data_w] = c766obus[data_w*3 +:data_w];
assign c766ibus[temp_w*4 +:temp_w] = v1918obus[temp_w*1 +:temp_w];
assign v1918ibus[data_w*1 +:data_w] = c766obus[data_w*4 +:data_w];
assign c766ibus[temp_w*5 +:temp_w] = v2014obus[temp_w*0 +:temp_w];
assign v2014ibus[data_w*0 +:data_w] = c766obus[data_w*5 +:data_w];
assign c767ibus[temp_w*0 +:temp_w] = v106obus[temp_w*2 +:temp_w];
assign v106ibus[data_w*2 +:data_w] = c767obus[data_w*0 +:data_w];
assign c767ibus[temp_w*1 +:temp_w] = v264obus[temp_w*4 +:temp_w];
assign v264ibus[data_w*4 +:data_w] = c767obus[data_w*1 +:data_w];
assign c767ibus[temp_w*2 +:temp_w] = v577obus[temp_w*2 +:temp_w];
assign v577ibus[data_w*2 +:data_w] = c767obus[data_w*2 +:data_w];
assign c767ibus[temp_w*3 +:temp_w] = v910obus[temp_w*4 +:temp_w];
assign v910ibus[data_w*4 +:data_w] = c767obus[data_w*3 +:data_w];
assign c767ibus[temp_w*4 +:temp_w] = v1919obus[temp_w*1 +:temp_w];
assign v1919ibus[data_w*1 +:data_w] = c767obus[data_w*4 +:data_w];
assign c767ibus[temp_w*5 +:temp_w] = v2015obus[temp_w*0 +:temp_w];
assign v2015ibus[data_w*0 +:data_w] = c767obus[data_w*5 +:data_w];
assign c768ibus[temp_w*0 +:temp_w] = v12obus[temp_w*1 +:temp_w];
assign v12ibus[data_w*1 +:data_w] = c768obus[data_w*0 +:data_w];
assign c768ibus[temp_w*1 +:temp_w] = v467obus[temp_w*2 +:temp_w];
assign v467ibus[data_w*2 +:data_w] = c768obus[data_w*1 +:data_w];
assign c768ibus[temp_w*2 +:temp_w] = v504obus[temp_w*3 +:temp_w];
assign v504ibus[data_w*3 +:data_w] = c768obus[data_w*2 +:data_w];
assign c768ibus[temp_w*3 +:temp_w] = v715obus[temp_w*3 +:temp_w];
assign v715ibus[data_w*3 +:data_w] = c768obus[data_w*3 +:data_w];
assign c768ibus[temp_w*4 +:temp_w] = v1107obus[temp_w*3 +:temp_w];
assign v1107ibus[data_w*3 +:data_w] = c768obus[data_w*4 +:data_w];
assign c768ibus[temp_w*5 +:temp_w] = v1920obus[temp_w*1 +:temp_w];
assign v1920ibus[data_w*1 +:data_w] = c768obus[data_w*5 +:data_w];
assign c768ibus[temp_w*6 +:temp_w] = v2016obus[temp_w*0 +:temp_w];
assign v2016ibus[data_w*0 +:data_w] = c768obus[data_w*6 +:data_w];
assign c769ibus[temp_w*0 +:temp_w] = v13obus[temp_w*1 +:temp_w];
assign v13ibus[data_w*1 +:data_w] = c769obus[data_w*0 +:data_w];
assign c769ibus[temp_w*1 +:temp_w] = v468obus[temp_w*2 +:temp_w];
assign v468ibus[data_w*2 +:data_w] = c769obus[data_w*1 +:data_w];
assign c769ibus[temp_w*2 +:temp_w] = v505obus[temp_w*3 +:temp_w];
assign v505ibus[data_w*3 +:data_w] = c769obus[data_w*2 +:data_w];
assign c769ibus[temp_w*3 +:temp_w] = v716obus[temp_w*3 +:temp_w];
assign v716ibus[data_w*3 +:data_w] = c769obus[data_w*3 +:data_w];
assign c769ibus[temp_w*4 +:temp_w] = v1108obus[temp_w*3 +:temp_w];
assign v1108ibus[data_w*3 +:data_w] = c769obus[data_w*4 +:data_w];
assign c769ibus[temp_w*5 +:temp_w] = v1921obus[temp_w*1 +:temp_w];
assign v1921ibus[data_w*1 +:data_w] = c769obus[data_w*5 +:data_w];
assign c769ibus[temp_w*6 +:temp_w] = v2017obus[temp_w*0 +:temp_w];
assign v2017ibus[data_w*0 +:data_w] = c769obus[data_w*6 +:data_w];
assign c770ibus[temp_w*0 +:temp_w] = v14obus[temp_w*1 +:temp_w];
assign v14ibus[data_w*1 +:data_w] = c770obus[data_w*0 +:data_w];
assign c770ibus[temp_w*1 +:temp_w] = v469obus[temp_w*2 +:temp_w];
assign v469ibus[data_w*2 +:data_w] = c770obus[data_w*1 +:data_w];
assign c770ibus[temp_w*2 +:temp_w] = v506obus[temp_w*3 +:temp_w];
assign v506ibus[data_w*3 +:data_w] = c770obus[data_w*2 +:data_w];
assign c770ibus[temp_w*3 +:temp_w] = v717obus[temp_w*3 +:temp_w];
assign v717ibus[data_w*3 +:data_w] = c770obus[data_w*3 +:data_w];
assign c770ibus[temp_w*4 +:temp_w] = v1109obus[temp_w*3 +:temp_w];
assign v1109ibus[data_w*3 +:data_w] = c770obus[data_w*4 +:data_w];
assign c770ibus[temp_w*5 +:temp_w] = v1922obus[temp_w*1 +:temp_w];
assign v1922ibus[data_w*1 +:data_w] = c770obus[data_w*5 +:data_w];
assign c770ibus[temp_w*6 +:temp_w] = v2018obus[temp_w*0 +:temp_w];
assign v2018ibus[data_w*0 +:data_w] = c770obus[data_w*6 +:data_w];
assign c771ibus[temp_w*0 +:temp_w] = v15obus[temp_w*1 +:temp_w];
assign v15ibus[data_w*1 +:data_w] = c771obus[data_w*0 +:data_w];
assign c771ibus[temp_w*1 +:temp_w] = v470obus[temp_w*2 +:temp_w];
assign v470ibus[data_w*2 +:data_w] = c771obus[data_w*1 +:data_w];
assign c771ibus[temp_w*2 +:temp_w] = v507obus[temp_w*3 +:temp_w];
assign v507ibus[data_w*3 +:data_w] = c771obus[data_w*2 +:data_w];
assign c771ibus[temp_w*3 +:temp_w] = v718obus[temp_w*3 +:temp_w];
assign v718ibus[data_w*3 +:data_w] = c771obus[data_w*3 +:data_w];
assign c771ibus[temp_w*4 +:temp_w] = v1110obus[temp_w*3 +:temp_w];
assign v1110ibus[data_w*3 +:data_w] = c771obus[data_w*4 +:data_w];
assign c771ibus[temp_w*5 +:temp_w] = v1923obus[temp_w*1 +:temp_w];
assign v1923ibus[data_w*1 +:data_w] = c771obus[data_w*5 +:data_w];
assign c771ibus[temp_w*6 +:temp_w] = v2019obus[temp_w*0 +:temp_w];
assign v2019ibus[data_w*0 +:data_w] = c771obus[data_w*6 +:data_w];
assign c772ibus[temp_w*0 +:temp_w] = v16obus[temp_w*1 +:temp_w];
assign v16ibus[data_w*1 +:data_w] = c772obus[data_w*0 +:data_w];
assign c772ibus[temp_w*1 +:temp_w] = v471obus[temp_w*2 +:temp_w];
assign v471ibus[data_w*2 +:data_w] = c772obus[data_w*1 +:data_w];
assign c772ibus[temp_w*2 +:temp_w] = v508obus[temp_w*3 +:temp_w];
assign v508ibus[data_w*3 +:data_w] = c772obus[data_w*2 +:data_w];
assign c772ibus[temp_w*3 +:temp_w] = v719obus[temp_w*3 +:temp_w];
assign v719ibus[data_w*3 +:data_w] = c772obus[data_w*3 +:data_w];
assign c772ibus[temp_w*4 +:temp_w] = v1111obus[temp_w*3 +:temp_w];
assign v1111ibus[data_w*3 +:data_w] = c772obus[data_w*4 +:data_w];
assign c772ibus[temp_w*5 +:temp_w] = v1924obus[temp_w*1 +:temp_w];
assign v1924ibus[data_w*1 +:data_w] = c772obus[data_w*5 +:data_w];
assign c772ibus[temp_w*6 +:temp_w] = v2020obus[temp_w*0 +:temp_w];
assign v2020ibus[data_w*0 +:data_w] = c772obus[data_w*6 +:data_w];
assign c773ibus[temp_w*0 +:temp_w] = v17obus[temp_w*1 +:temp_w];
assign v17ibus[data_w*1 +:data_w] = c773obus[data_w*0 +:data_w];
assign c773ibus[temp_w*1 +:temp_w] = v472obus[temp_w*2 +:temp_w];
assign v472ibus[data_w*2 +:data_w] = c773obus[data_w*1 +:data_w];
assign c773ibus[temp_w*2 +:temp_w] = v509obus[temp_w*3 +:temp_w];
assign v509ibus[data_w*3 +:data_w] = c773obus[data_w*2 +:data_w];
assign c773ibus[temp_w*3 +:temp_w] = v720obus[temp_w*3 +:temp_w];
assign v720ibus[data_w*3 +:data_w] = c773obus[data_w*3 +:data_w];
assign c773ibus[temp_w*4 +:temp_w] = v1112obus[temp_w*3 +:temp_w];
assign v1112ibus[data_w*3 +:data_w] = c773obus[data_w*4 +:data_w];
assign c773ibus[temp_w*5 +:temp_w] = v1925obus[temp_w*1 +:temp_w];
assign v1925ibus[data_w*1 +:data_w] = c773obus[data_w*5 +:data_w];
assign c773ibus[temp_w*6 +:temp_w] = v2021obus[temp_w*0 +:temp_w];
assign v2021ibus[data_w*0 +:data_w] = c773obus[data_w*6 +:data_w];
assign c774ibus[temp_w*0 +:temp_w] = v18obus[temp_w*1 +:temp_w];
assign v18ibus[data_w*1 +:data_w] = c774obus[data_w*0 +:data_w];
assign c774ibus[temp_w*1 +:temp_w] = v473obus[temp_w*2 +:temp_w];
assign v473ibus[data_w*2 +:data_w] = c774obus[data_w*1 +:data_w];
assign c774ibus[temp_w*2 +:temp_w] = v510obus[temp_w*3 +:temp_w];
assign v510ibus[data_w*3 +:data_w] = c774obus[data_w*2 +:data_w];
assign c774ibus[temp_w*3 +:temp_w] = v721obus[temp_w*3 +:temp_w];
assign v721ibus[data_w*3 +:data_w] = c774obus[data_w*3 +:data_w];
assign c774ibus[temp_w*4 +:temp_w] = v1113obus[temp_w*3 +:temp_w];
assign v1113ibus[data_w*3 +:data_w] = c774obus[data_w*4 +:data_w];
assign c774ibus[temp_w*5 +:temp_w] = v1926obus[temp_w*1 +:temp_w];
assign v1926ibus[data_w*1 +:data_w] = c774obus[data_w*5 +:data_w];
assign c774ibus[temp_w*6 +:temp_w] = v2022obus[temp_w*0 +:temp_w];
assign v2022ibus[data_w*0 +:data_w] = c774obus[data_w*6 +:data_w];
assign c775ibus[temp_w*0 +:temp_w] = v19obus[temp_w*1 +:temp_w];
assign v19ibus[data_w*1 +:data_w] = c775obus[data_w*0 +:data_w];
assign c775ibus[temp_w*1 +:temp_w] = v474obus[temp_w*2 +:temp_w];
assign v474ibus[data_w*2 +:data_w] = c775obus[data_w*1 +:data_w];
assign c775ibus[temp_w*2 +:temp_w] = v511obus[temp_w*3 +:temp_w];
assign v511ibus[data_w*3 +:data_w] = c775obus[data_w*2 +:data_w];
assign c775ibus[temp_w*3 +:temp_w] = v722obus[temp_w*3 +:temp_w];
assign v722ibus[data_w*3 +:data_w] = c775obus[data_w*3 +:data_w];
assign c775ibus[temp_w*4 +:temp_w] = v1114obus[temp_w*3 +:temp_w];
assign v1114ibus[data_w*3 +:data_w] = c775obus[data_w*4 +:data_w];
assign c775ibus[temp_w*5 +:temp_w] = v1927obus[temp_w*1 +:temp_w];
assign v1927ibus[data_w*1 +:data_w] = c775obus[data_w*5 +:data_w];
assign c775ibus[temp_w*6 +:temp_w] = v2023obus[temp_w*0 +:temp_w];
assign v2023ibus[data_w*0 +:data_w] = c775obus[data_w*6 +:data_w];
assign c776ibus[temp_w*0 +:temp_w] = v20obus[temp_w*1 +:temp_w];
assign v20ibus[data_w*1 +:data_w] = c776obus[data_w*0 +:data_w];
assign c776ibus[temp_w*1 +:temp_w] = v475obus[temp_w*2 +:temp_w];
assign v475ibus[data_w*2 +:data_w] = c776obus[data_w*1 +:data_w];
assign c776ibus[temp_w*2 +:temp_w] = v512obus[temp_w*3 +:temp_w];
assign v512ibus[data_w*3 +:data_w] = c776obus[data_w*2 +:data_w];
assign c776ibus[temp_w*3 +:temp_w] = v723obus[temp_w*3 +:temp_w];
assign v723ibus[data_w*3 +:data_w] = c776obus[data_w*3 +:data_w];
assign c776ibus[temp_w*4 +:temp_w] = v1115obus[temp_w*3 +:temp_w];
assign v1115ibus[data_w*3 +:data_w] = c776obus[data_w*4 +:data_w];
assign c776ibus[temp_w*5 +:temp_w] = v1928obus[temp_w*1 +:temp_w];
assign v1928ibus[data_w*1 +:data_w] = c776obus[data_w*5 +:data_w];
assign c776ibus[temp_w*6 +:temp_w] = v2024obus[temp_w*0 +:temp_w];
assign v2024ibus[data_w*0 +:data_w] = c776obus[data_w*6 +:data_w];
assign c777ibus[temp_w*0 +:temp_w] = v21obus[temp_w*1 +:temp_w];
assign v21ibus[data_w*1 +:data_w] = c777obus[data_w*0 +:data_w];
assign c777ibus[temp_w*1 +:temp_w] = v476obus[temp_w*2 +:temp_w];
assign v476ibus[data_w*2 +:data_w] = c777obus[data_w*1 +:data_w];
assign c777ibus[temp_w*2 +:temp_w] = v513obus[temp_w*3 +:temp_w];
assign v513ibus[data_w*3 +:data_w] = c777obus[data_w*2 +:data_w];
assign c777ibus[temp_w*3 +:temp_w] = v724obus[temp_w*3 +:temp_w];
assign v724ibus[data_w*3 +:data_w] = c777obus[data_w*3 +:data_w];
assign c777ibus[temp_w*4 +:temp_w] = v1116obus[temp_w*3 +:temp_w];
assign v1116ibus[data_w*3 +:data_w] = c777obus[data_w*4 +:data_w];
assign c777ibus[temp_w*5 +:temp_w] = v1929obus[temp_w*1 +:temp_w];
assign v1929ibus[data_w*1 +:data_w] = c777obus[data_w*5 +:data_w];
assign c777ibus[temp_w*6 +:temp_w] = v2025obus[temp_w*0 +:temp_w];
assign v2025ibus[data_w*0 +:data_w] = c777obus[data_w*6 +:data_w];
assign c778ibus[temp_w*0 +:temp_w] = v22obus[temp_w*1 +:temp_w];
assign v22ibus[data_w*1 +:data_w] = c778obus[data_w*0 +:data_w];
assign c778ibus[temp_w*1 +:temp_w] = v477obus[temp_w*2 +:temp_w];
assign v477ibus[data_w*2 +:data_w] = c778obus[data_w*1 +:data_w];
assign c778ibus[temp_w*2 +:temp_w] = v514obus[temp_w*3 +:temp_w];
assign v514ibus[data_w*3 +:data_w] = c778obus[data_w*2 +:data_w];
assign c778ibus[temp_w*3 +:temp_w] = v725obus[temp_w*3 +:temp_w];
assign v725ibus[data_w*3 +:data_w] = c778obus[data_w*3 +:data_w];
assign c778ibus[temp_w*4 +:temp_w] = v1117obus[temp_w*3 +:temp_w];
assign v1117ibus[data_w*3 +:data_w] = c778obus[data_w*4 +:data_w];
assign c778ibus[temp_w*5 +:temp_w] = v1930obus[temp_w*1 +:temp_w];
assign v1930ibus[data_w*1 +:data_w] = c778obus[data_w*5 +:data_w];
assign c778ibus[temp_w*6 +:temp_w] = v2026obus[temp_w*0 +:temp_w];
assign v2026ibus[data_w*0 +:data_w] = c778obus[data_w*6 +:data_w];
assign c779ibus[temp_w*0 +:temp_w] = v23obus[temp_w*1 +:temp_w];
assign v23ibus[data_w*1 +:data_w] = c779obus[data_w*0 +:data_w];
assign c779ibus[temp_w*1 +:temp_w] = v478obus[temp_w*2 +:temp_w];
assign v478ibus[data_w*2 +:data_w] = c779obus[data_w*1 +:data_w];
assign c779ibus[temp_w*2 +:temp_w] = v515obus[temp_w*3 +:temp_w];
assign v515ibus[data_w*3 +:data_w] = c779obus[data_w*2 +:data_w];
assign c779ibus[temp_w*3 +:temp_w] = v726obus[temp_w*3 +:temp_w];
assign v726ibus[data_w*3 +:data_w] = c779obus[data_w*3 +:data_w];
assign c779ibus[temp_w*4 +:temp_w] = v1118obus[temp_w*3 +:temp_w];
assign v1118ibus[data_w*3 +:data_w] = c779obus[data_w*4 +:data_w];
assign c779ibus[temp_w*5 +:temp_w] = v1931obus[temp_w*1 +:temp_w];
assign v1931ibus[data_w*1 +:data_w] = c779obus[data_w*5 +:data_w];
assign c779ibus[temp_w*6 +:temp_w] = v2027obus[temp_w*0 +:temp_w];
assign v2027ibus[data_w*0 +:data_w] = c779obus[data_w*6 +:data_w];
assign c780ibus[temp_w*0 +:temp_w] = v24obus[temp_w*1 +:temp_w];
assign v24ibus[data_w*1 +:data_w] = c780obus[data_w*0 +:data_w];
assign c780ibus[temp_w*1 +:temp_w] = v479obus[temp_w*2 +:temp_w];
assign v479ibus[data_w*2 +:data_w] = c780obus[data_w*1 +:data_w];
assign c780ibus[temp_w*2 +:temp_w] = v516obus[temp_w*3 +:temp_w];
assign v516ibus[data_w*3 +:data_w] = c780obus[data_w*2 +:data_w];
assign c780ibus[temp_w*3 +:temp_w] = v727obus[temp_w*3 +:temp_w];
assign v727ibus[data_w*3 +:data_w] = c780obus[data_w*3 +:data_w];
assign c780ibus[temp_w*4 +:temp_w] = v1119obus[temp_w*3 +:temp_w];
assign v1119ibus[data_w*3 +:data_w] = c780obus[data_w*4 +:data_w];
assign c780ibus[temp_w*5 +:temp_w] = v1932obus[temp_w*1 +:temp_w];
assign v1932ibus[data_w*1 +:data_w] = c780obus[data_w*5 +:data_w];
assign c780ibus[temp_w*6 +:temp_w] = v2028obus[temp_w*0 +:temp_w];
assign v2028ibus[data_w*0 +:data_w] = c780obus[data_w*6 +:data_w];
assign c781ibus[temp_w*0 +:temp_w] = v25obus[temp_w*1 +:temp_w];
assign v25ibus[data_w*1 +:data_w] = c781obus[data_w*0 +:data_w];
assign c781ibus[temp_w*1 +:temp_w] = v384obus[temp_w*2 +:temp_w];
assign v384ibus[data_w*2 +:data_w] = c781obus[data_w*1 +:data_w];
assign c781ibus[temp_w*2 +:temp_w] = v517obus[temp_w*3 +:temp_w];
assign v517ibus[data_w*3 +:data_w] = c781obus[data_w*2 +:data_w];
assign c781ibus[temp_w*3 +:temp_w] = v728obus[temp_w*3 +:temp_w];
assign v728ibus[data_w*3 +:data_w] = c781obus[data_w*3 +:data_w];
assign c781ibus[temp_w*4 +:temp_w] = v1120obus[temp_w*3 +:temp_w];
assign v1120ibus[data_w*3 +:data_w] = c781obus[data_w*4 +:data_w];
assign c781ibus[temp_w*5 +:temp_w] = v1933obus[temp_w*1 +:temp_w];
assign v1933ibus[data_w*1 +:data_w] = c781obus[data_w*5 +:data_w];
assign c781ibus[temp_w*6 +:temp_w] = v2029obus[temp_w*0 +:temp_w];
assign v2029ibus[data_w*0 +:data_w] = c781obus[data_w*6 +:data_w];
assign c782ibus[temp_w*0 +:temp_w] = v26obus[temp_w*1 +:temp_w];
assign v26ibus[data_w*1 +:data_w] = c782obus[data_w*0 +:data_w];
assign c782ibus[temp_w*1 +:temp_w] = v385obus[temp_w*2 +:temp_w];
assign v385ibus[data_w*2 +:data_w] = c782obus[data_w*1 +:data_w];
assign c782ibus[temp_w*2 +:temp_w] = v518obus[temp_w*3 +:temp_w];
assign v518ibus[data_w*3 +:data_w] = c782obus[data_w*2 +:data_w];
assign c782ibus[temp_w*3 +:temp_w] = v729obus[temp_w*3 +:temp_w];
assign v729ibus[data_w*3 +:data_w] = c782obus[data_w*3 +:data_w];
assign c782ibus[temp_w*4 +:temp_w] = v1121obus[temp_w*3 +:temp_w];
assign v1121ibus[data_w*3 +:data_w] = c782obus[data_w*4 +:data_w];
assign c782ibus[temp_w*5 +:temp_w] = v1934obus[temp_w*1 +:temp_w];
assign v1934ibus[data_w*1 +:data_w] = c782obus[data_w*5 +:data_w];
assign c782ibus[temp_w*6 +:temp_w] = v2030obus[temp_w*0 +:temp_w];
assign v2030ibus[data_w*0 +:data_w] = c782obus[data_w*6 +:data_w];
assign c783ibus[temp_w*0 +:temp_w] = v27obus[temp_w*1 +:temp_w];
assign v27ibus[data_w*1 +:data_w] = c783obus[data_w*0 +:data_w];
assign c783ibus[temp_w*1 +:temp_w] = v386obus[temp_w*2 +:temp_w];
assign v386ibus[data_w*2 +:data_w] = c783obus[data_w*1 +:data_w];
assign c783ibus[temp_w*2 +:temp_w] = v519obus[temp_w*3 +:temp_w];
assign v519ibus[data_w*3 +:data_w] = c783obus[data_w*2 +:data_w];
assign c783ibus[temp_w*3 +:temp_w] = v730obus[temp_w*3 +:temp_w];
assign v730ibus[data_w*3 +:data_w] = c783obus[data_w*3 +:data_w];
assign c783ibus[temp_w*4 +:temp_w] = v1122obus[temp_w*3 +:temp_w];
assign v1122ibus[data_w*3 +:data_w] = c783obus[data_w*4 +:data_w];
assign c783ibus[temp_w*5 +:temp_w] = v1935obus[temp_w*1 +:temp_w];
assign v1935ibus[data_w*1 +:data_w] = c783obus[data_w*5 +:data_w];
assign c783ibus[temp_w*6 +:temp_w] = v2031obus[temp_w*0 +:temp_w];
assign v2031ibus[data_w*0 +:data_w] = c783obus[data_w*6 +:data_w];
assign c784ibus[temp_w*0 +:temp_w] = v28obus[temp_w*1 +:temp_w];
assign v28ibus[data_w*1 +:data_w] = c784obus[data_w*0 +:data_w];
assign c784ibus[temp_w*1 +:temp_w] = v387obus[temp_w*2 +:temp_w];
assign v387ibus[data_w*2 +:data_w] = c784obus[data_w*1 +:data_w];
assign c784ibus[temp_w*2 +:temp_w] = v520obus[temp_w*3 +:temp_w];
assign v520ibus[data_w*3 +:data_w] = c784obus[data_w*2 +:data_w];
assign c784ibus[temp_w*3 +:temp_w] = v731obus[temp_w*3 +:temp_w];
assign v731ibus[data_w*3 +:data_w] = c784obus[data_w*3 +:data_w];
assign c784ibus[temp_w*4 +:temp_w] = v1123obus[temp_w*3 +:temp_w];
assign v1123ibus[data_w*3 +:data_w] = c784obus[data_w*4 +:data_w];
assign c784ibus[temp_w*5 +:temp_w] = v1936obus[temp_w*1 +:temp_w];
assign v1936ibus[data_w*1 +:data_w] = c784obus[data_w*5 +:data_w];
assign c784ibus[temp_w*6 +:temp_w] = v2032obus[temp_w*0 +:temp_w];
assign v2032ibus[data_w*0 +:data_w] = c784obus[data_w*6 +:data_w];
assign c785ibus[temp_w*0 +:temp_w] = v29obus[temp_w*1 +:temp_w];
assign v29ibus[data_w*1 +:data_w] = c785obus[data_w*0 +:data_w];
assign c785ibus[temp_w*1 +:temp_w] = v388obus[temp_w*2 +:temp_w];
assign v388ibus[data_w*2 +:data_w] = c785obus[data_w*1 +:data_w];
assign c785ibus[temp_w*2 +:temp_w] = v521obus[temp_w*3 +:temp_w];
assign v521ibus[data_w*3 +:data_w] = c785obus[data_w*2 +:data_w];
assign c785ibus[temp_w*3 +:temp_w] = v732obus[temp_w*3 +:temp_w];
assign v732ibus[data_w*3 +:data_w] = c785obus[data_w*3 +:data_w];
assign c785ibus[temp_w*4 +:temp_w] = v1124obus[temp_w*3 +:temp_w];
assign v1124ibus[data_w*3 +:data_w] = c785obus[data_w*4 +:data_w];
assign c785ibus[temp_w*5 +:temp_w] = v1937obus[temp_w*1 +:temp_w];
assign v1937ibus[data_w*1 +:data_w] = c785obus[data_w*5 +:data_w];
assign c785ibus[temp_w*6 +:temp_w] = v2033obus[temp_w*0 +:temp_w];
assign v2033ibus[data_w*0 +:data_w] = c785obus[data_w*6 +:data_w];
assign c786ibus[temp_w*0 +:temp_w] = v30obus[temp_w*1 +:temp_w];
assign v30ibus[data_w*1 +:data_w] = c786obus[data_w*0 +:data_w];
assign c786ibus[temp_w*1 +:temp_w] = v389obus[temp_w*2 +:temp_w];
assign v389ibus[data_w*2 +:data_w] = c786obus[data_w*1 +:data_w];
assign c786ibus[temp_w*2 +:temp_w] = v522obus[temp_w*3 +:temp_w];
assign v522ibus[data_w*3 +:data_w] = c786obus[data_w*2 +:data_w];
assign c786ibus[temp_w*3 +:temp_w] = v733obus[temp_w*3 +:temp_w];
assign v733ibus[data_w*3 +:data_w] = c786obus[data_w*3 +:data_w];
assign c786ibus[temp_w*4 +:temp_w] = v1125obus[temp_w*3 +:temp_w];
assign v1125ibus[data_w*3 +:data_w] = c786obus[data_w*4 +:data_w];
assign c786ibus[temp_w*5 +:temp_w] = v1938obus[temp_w*1 +:temp_w];
assign v1938ibus[data_w*1 +:data_w] = c786obus[data_w*5 +:data_w];
assign c786ibus[temp_w*6 +:temp_w] = v2034obus[temp_w*0 +:temp_w];
assign v2034ibus[data_w*0 +:data_w] = c786obus[data_w*6 +:data_w];
assign c787ibus[temp_w*0 +:temp_w] = v31obus[temp_w*1 +:temp_w];
assign v31ibus[data_w*1 +:data_w] = c787obus[data_w*0 +:data_w];
assign c787ibus[temp_w*1 +:temp_w] = v390obus[temp_w*2 +:temp_w];
assign v390ibus[data_w*2 +:data_w] = c787obus[data_w*1 +:data_w];
assign c787ibus[temp_w*2 +:temp_w] = v523obus[temp_w*3 +:temp_w];
assign v523ibus[data_w*3 +:data_w] = c787obus[data_w*2 +:data_w];
assign c787ibus[temp_w*3 +:temp_w] = v734obus[temp_w*3 +:temp_w];
assign v734ibus[data_w*3 +:data_w] = c787obus[data_w*3 +:data_w];
assign c787ibus[temp_w*4 +:temp_w] = v1126obus[temp_w*3 +:temp_w];
assign v1126ibus[data_w*3 +:data_w] = c787obus[data_w*4 +:data_w];
assign c787ibus[temp_w*5 +:temp_w] = v1939obus[temp_w*1 +:temp_w];
assign v1939ibus[data_w*1 +:data_w] = c787obus[data_w*5 +:data_w];
assign c787ibus[temp_w*6 +:temp_w] = v2035obus[temp_w*0 +:temp_w];
assign v2035ibus[data_w*0 +:data_w] = c787obus[data_w*6 +:data_w];
assign c788ibus[temp_w*0 +:temp_w] = v32obus[temp_w*1 +:temp_w];
assign v32ibus[data_w*1 +:data_w] = c788obus[data_w*0 +:data_w];
assign c788ibus[temp_w*1 +:temp_w] = v391obus[temp_w*2 +:temp_w];
assign v391ibus[data_w*2 +:data_w] = c788obus[data_w*1 +:data_w];
assign c788ibus[temp_w*2 +:temp_w] = v524obus[temp_w*3 +:temp_w];
assign v524ibus[data_w*3 +:data_w] = c788obus[data_w*2 +:data_w];
assign c788ibus[temp_w*3 +:temp_w] = v735obus[temp_w*3 +:temp_w];
assign v735ibus[data_w*3 +:data_w] = c788obus[data_w*3 +:data_w];
assign c788ibus[temp_w*4 +:temp_w] = v1127obus[temp_w*3 +:temp_w];
assign v1127ibus[data_w*3 +:data_w] = c788obus[data_w*4 +:data_w];
assign c788ibus[temp_w*5 +:temp_w] = v1940obus[temp_w*1 +:temp_w];
assign v1940ibus[data_w*1 +:data_w] = c788obus[data_w*5 +:data_w];
assign c788ibus[temp_w*6 +:temp_w] = v2036obus[temp_w*0 +:temp_w];
assign v2036ibus[data_w*0 +:data_w] = c788obus[data_w*6 +:data_w];
assign c789ibus[temp_w*0 +:temp_w] = v33obus[temp_w*1 +:temp_w];
assign v33ibus[data_w*1 +:data_w] = c789obus[data_w*0 +:data_w];
assign c789ibus[temp_w*1 +:temp_w] = v392obus[temp_w*2 +:temp_w];
assign v392ibus[data_w*2 +:data_w] = c789obus[data_w*1 +:data_w];
assign c789ibus[temp_w*2 +:temp_w] = v525obus[temp_w*3 +:temp_w];
assign v525ibus[data_w*3 +:data_w] = c789obus[data_w*2 +:data_w];
assign c789ibus[temp_w*3 +:temp_w] = v736obus[temp_w*3 +:temp_w];
assign v736ibus[data_w*3 +:data_w] = c789obus[data_w*3 +:data_w];
assign c789ibus[temp_w*4 +:temp_w] = v1128obus[temp_w*3 +:temp_w];
assign v1128ibus[data_w*3 +:data_w] = c789obus[data_w*4 +:data_w];
assign c789ibus[temp_w*5 +:temp_w] = v1941obus[temp_w*1 +:temp_w];
assign v1941ibus[data_w*1 +:data_w] = c789obus[data_w*5 +:data_w];
assign c789ibus[temp_w*6 +:temp_w] = v2037obus[temp_w*0 +:temp_w];
assign v2037ibus[data_w*0 +:data_w] = c789obus[data_w*6 +:data_w];
assign c790ibus[temp_w*0 +:temp_w] = v34obus[temp_w*1 +:temp_w];
assign v34ibus[data_w*1 +:data_w] = c790obus[data_w*0 +:data_w];
assign c790ibus[temp_w*1 +:temp_w] = v393obus[temp_w*2 +:temp_w];
assign v393ibus[data_w*2 +:data_w] = c790obus[data_w*1 +:data_w];
assign c790ibus[temp_w*2 +:temp_w] = v526obus[temp_w*3 +:temp_w];
assign v526ibus[data_w*3 +:data_w] = c790obus[data_w*2 +:data_w];
assign c790ibus[temp_w*3 +:temp_w] = v737obus[temp_w*3 +:temp_w];
assign v737ibus[data_w*3 +:data_w] = c790obus[data_w*3 +:data_w];
assign c790ibus[temp_w*4 +:temp_w] = v1129obus[temp_w*3 +:temp_w];
assign v1129ibus[data_w*3 +:data_w] = c790obus[data_w*4 +:data_w];
assign c790ibus[temp_w*5 +:temp_w] = v1942obus[temp_w*1 +:temp_w];
assign v1942ibus[data_w*1 +:data_w] = c790obus[data_w*5 +:data_w];
assign c790ibus[temp_w*6 +:temp_w] = v2038obus[temp_w*0 +:temp_w];
assign v2038ibus[data_w*0 +:data_w] = c790obus[data_w*6 +:data_w];
assign c791ibus[temp_w*0 +:temp_w] = v35obus[temp_w*1 +:temp_w];
assign v35ibus[data_w*1 +:data_w] = c791obus[data_w*0 +:data_w];
assign c791ibus[temp_w*1 +:temp_w] = v394obus[temp_w*2 +:temp_w];
assign v394ibus[data_w*2 +:data_w] = c791obus[data_w*1 +:data_w];
assign c791ibus[temp_w*2 +:temp_w] = v527obus[temp_w*3 +:temp_w];
assign v527ibus[data_w*3 +:data_w] = c791obus[data_w*2 +:data_w];
assign c791ibus[temp_w*3 +:temp_w] = v738obus[temp_w*3 +:temp_w];
assign v738ibus[data_w*3 +:data_w] = c791obus[data_w*3 +:data_w];
assign c791ibus[temp_w*4 +:temp_w] = v1130obus[temp_w*3 +:temp_w];
assign v1130ibus[data_w*3 +:data_w] = c791obus[data_w*4 +:data_w];
assign c791ibus[temp_w*5 +:temp_w] = v1943obus[temp_w*1 +:temp_w];
assign v1943ibus[data_w*1 +:data_w] = c791obus[data_w*5 +:data_w];
assign c791ibus[temp_w*6 +:temp_w] = v2039obus[temp_w*0 +:temp_w];
assign v2039ibus[data_w*0 +:data_w] = c791obus[data_w*6 +:data_w];
assign c792ibus[temp_w*0 +:temp_w] = v36obus[temp_w*1 +:temp_w];
assign v36ibus[data_w*1 +:data_w] = c792obus[data_w*0 +:data_w];
assign c792ibus[temp_w*1 +:temp_w] = v395obus[temp_w*2 +:temp_w];
assign v395ibus[data_w*2 +:data_w] = c792obus[data_w*1 +:data_w];
assign c792ibus[temp_w*2 +:temp_w] = v528obus[temp_w*3 +:temp_w];
assign v528ibus[data_w*3 +:data_w] = c792obus[data_w*2 +:data_w];
assign c792ibus[temp_w*3 +:temp_w] = v739obus[temp_w*3 +:temp_w];
assign v739ibus[data_w*3 +:data_w] = c792obus[data_w*3 +:data_w];
assign c792ibus[temp_w*4 +:temp_w] = v1131obus[temp_w*3 +:temp_w];
assign v1131ibus[data_w*3 +:data_w] = c792obus[data_w*4 +:data_w];
assign c792ibus[temp_w*5 +:temp_w] = v1944obus[temp_w*1 +:temp_w];
assign v1944ibus[data_w*1 +:data_w] = c792obus[data_w*5 +:data_w];
assign c792ibus[temp_w*6 +:temp_w] = v2040obus[temp_w*0 +:temp_w];
assign v2040ibus[data_w*0 +:data_w] = c792obus[data_w*6 +:data_w];
assign c793ibus[temp_w*0 +:temp_w] = v37obus[temp_w*1 +:temp_w];
assign v37ibus[data_w*1 +:data_w] = c793obus[data_w*0 +:data_w];
assign c793ibus[temp_w*1 +:temp_w] = v396obus[temp_w*2 +:temp_w];
assign v396ibus[data_w*2 +:data_w] = c793obus[data_w*1 +:data_w];
assign c793ibus[temp_w*2 +:temp_w] = v529obus[temp_w*3 +:temp_w];
assign v529ibus[data_w*3 +:data_w] = c793obus[data_w*2 +:data_w];
assign c793ibus[temp_w*3 +:temp_w] = v740obus[temp_w*3 +:temp_w];
assign v740ibus[data_w*3 +:data_w] = c793obus[data_w*3 +:data_w];
assign c793ibus[temp_w*4 +:temp_w] = v1132obus[temp_w*3 +:temp_w];
assign v1132ibus[data_w*3 +:data_w] = c793obus[data_w*4 +:data_w];
assign c793ibus[temp_w*5 +:temp_w] = v1945obus[temp_w*1 +:temp_w];
assign v1945ibus[data_w*1 +:data_w] = c793obus[data_w*5 +:data_w];
assign c793ibus[temp_w*6 +:temp_w] = v2041obus[temp_w*0 +:temp_w];
assign v2041ibus[data_w*0 +:data_w] = c793obus[data_w*6 +:data_w];
assign c794ibus[temp_w*0 +:temp_w] = v38obus[temp_w*1 +:temp_w];
assign v38ibus[data_w*1 +:data_w] = c794obus[data_w*0 +:data_w];
assign c794ibus[temp_w*1 +:temp_w] = v397obus[temp_w*2 +:temp_w];
assign v397ibus[data_w*2 +:data_w] = c794obus[data_w*1 +:data_w];
assign c794ibus[temp_w*2 +:temp_w] = v530obus[temp_w*3 +:temp_w];
assign v530ibus[data_w*3 +:data_w] = c794obus[data_w*2 +:data_w];
assign c794ibus[temp_w*3 +:temp_w] = v741obus[temp_w*3 +:temp_w];
assign v741ibus[data_w*3 +:data_w] = c794obus[data_w*3 +:data_w];
assign c794ibus[temp_w*4 +:temp_w] = v1133obus[temp_w*3 +:temp_w];
assign v1133ibus[data_w*3 +:data_w] = c794obus[data_w*4 +:data_w];
assign c794ibus[temp_w*5 +:temp_w] = v1946obus[temp_w*1 +:temp_w];
assign v1946ibus[data_w*1 +:data_w] = c794obus[data_w*5 +:data_w];
assign c794ibus[temp_w*6 +:temp_w] = v2042obus[temp_w*0 +:temp_w];
assign v2042ibus[data_w*0 +:data_w] = c794obus[data_w*6 +:data_w];
assign c795ibus[temp_w*0 +:temp_w] = v39obus[temp_w*1 +:temp_w];
assign v39ibus[data_w*1 +:data_w] = c795obus[data_w*0 +:data_w];
assign c795ibus[temp_w*1 +:temp_w] = v398obus[temp_w*2 +:temp_w];
assign v398ibus[data_w*2 +:data_w] = c795obus[data_w*1 +:data_w];
assign c795ibus[temp_w*2 +:temp_w] = v531obus[temp_w*3 +:temp_w];
assign v531ibus[data_w*3 +:data_w] = c795obus[data_w*2 +:data_w];
assign c795ibus[temp_w*3 +:temp_w] = v742obus[temp_w*3 +:temp_w];
assign v742ibus[data_w*3 +:data_w] = c795obus[data_w*3 +:data_w];
assign c795ibus[temp_w*4 +:temp_w] = v1134obus[temp_w*3 +:temp_w];
assign v1134ibus[data_w*3 +:data_w] = c795obus[data_w*4 +:data_w];
assign c795ibus[temp_w*5 +:temp_w] = v1947obus[temp_w*1 +:temp_w];
assign v1947ibus[data_w*1 +:data_w] = c795obus[data_w*5 +:data_w];
assign c795ibus[temp_w*6 +:temp_w] = v2043obus[temp_w*0 +:temp_w];
assign v2043ibus[data_w*0 +:data_w] = c795obus[data_w*6 +:data_w];
assign c796ibus[temp_w*0 +:temp_w] = v40obus[temp_w*1 +:temp_w];
assign v40ibus[data_w*1 +:data_w] = c796obus[data_w*0 +:data_w];
assign c796ibus[temp_w*1 +:temp_w] = v399obus[temp_w*2 +:temp_w];
assign v399ibus[data_w*2 +:data_w] = c796obus[data_w*1 +:data_w];
assign c796ibus[temp_w*2 +:temp_w] = v532obus[temp_w*3 +:temp_w];
assign v532ibus[data_w*3 +:data_w] = c796obus[data_w*2 +:data_w];
assign c796ibus[temp_w*3 +:temp_w] = v743obus[temp_w*3 +:temp_w];
assign v743ibus[data_w*3 +:data_w] = c796obus[data_w*3 +:data_w];
assign c796ibus[temp_w*4 +:temp_w] = v1135obus[temp_w*3 +:temp_w];
assign v1135ibus[data_w*3 +:data_w] = c796obus[data_w*4 +:data_w];
assign c796ibus[temp_w*5 +:temp_w] = v1948obus[temp_w*1 +:temp_w];
assign v1948ibus[data_w*1 +:data_w] = c796obus[data_w*5 +:data_w];
assign c796ibus[temp_w*6 +:temp_w] = v2044obus[temp_w*0 +:temp_w];
assign v2044ibus[data_w*0 +:data_w] = c796obus[data_w*6 +:data_w];
assign c797ibus[temp_w*0 +:temp_w] = v41obus[temp_w*1 +:temp_w];
assign v41ibus[data_w*1 +:data_w] = c797obus[data_w*0 +:data_w];
assign c797ibus[temp_w*1 +:temp_w] = v400obus[temp_w*2 +:temp_w];
assign v400ibus[data_w*2 +:data_w] = c797obus[data_w*1 +:data_w];
assign c797ibus[temp_w*2 +:temp_w] = v533obus[temp_w*3 +:temp_w];
assign v533ibus[data_w*3 +:data_w] = c797obus[data_w*2 +:data_w];
assign c797ibus[temp_w*3 +:temp_w] = v744obus[temp_w*3 +:temp_w];
assign v744ibus[data_w*3 +:data_w] = c797obus[data_w*3 +:data_w];
assign c797ibus[temp_w*4 +:temp_w] = v1136obus[temp_w*3 +:temp_w];
assign v1136ibus[data_w*3 +:data_w] = c797obus[data_w*4 +:data_w];
assign c797ibus[temp_w*5 +:temp_w] = v1949obus[temp_w*1 +:temp_w];
assign v1949ibus[data_w*1 +:data_w] = c797obus[data_w*5 +:data_w];
assign c797ibus[temp_w*6 +:temp_w] = v2045obus[temp_w*0 +:temp_w];
assign v2045ibus[data_w*0 +:data_w] = c797obus[data_w*6 +:data_w];
assign c798ibus[temp_w*0 +:temp_w] = v42obus[temp_w*1 +:temp_w];
assign v42ibus[data_w*1 +:data_w] = c798obus[data_w*0 +:data_w];
assign c798ibus[temp_w*1 +:temp_w] = v401obus[temp_w*2 +:temp_w];
assign v401ibus[data_w*2 +:data_w] = c798obus[data_w*1 +:data_w];
assign c798ibus[temp_w*2 +:temp_w] = v534obus[temp_w*3 +:temp_w];
assign v534ibus[data_w*3 +:data_w] = c798obus[data_w*2 +:data_w];
assign c798ibus[temp_w*3 +:temp_w] = v745obus[temp_w*3 +:temp_w];
assign v745ibus[data_w*3 +:data_w] = c798obus[data_w*3 +:data_w];
assign c798ibus[temp_w*4 +:temp_w] = v1137obus[temp_w*3 +:temp_w];
assign v1137ibus[data_w*3 +:data_w] = c798obus[data_w*4 +:data_w];
assign c798ibus[temp_w*5 +:temp_w] = v1950obus[temp_w*1 +:temp_w];
assign v1950ibus[data_w*1 +:data_w] = c798obus[data_w*5 +:data_w];
assign c798ibus[temp_w*6 +:temp_w] = v2046obus[temp_w*0 +:temp_w];
assign v2046ibus[data_w*0 +:data_w] = c798obus[data_w*6 +:data_w];
assign c799ibus[temp_w*0 +:temp_w] = v43obus[temp_w*1 +:temp_w];
assign v43ibus[data_w*1 +:data_w] = c799obus[data_w*0 +:data_w];
assign c799ibus[temp_w*1 +:temp_w] = v402obus[temp_w*2 +:temp_w];
assign v402ibus[data_w*2 +:data_w] = c799obus[data_w*1 +:data_w];
assign c799ibus[temp_w*2 +:temp_w] = v535obus[temp_w*3 +:temp_w];
assign v535ibus[data_w*3 +:data_w] = c799obus[data_w*2 +:data_w];
assign c799ibus[temp_w*3 +:temp_w] = v746obus[temp_w*3 +:temp_w];
assign v746ibus[data_w*3 +:data_w] = c799obus[data_w*3 +:data_w];
assign c799ibus[temp_w*4 +:temp_w] = v1138obus[temp_w*3 +:temp_w];
assign v1138ibus[data_w*3 +:data_w] = c799obus[data_w*4 +:data_w];
assign c799ibus[temp_w*5 +:temp_w] = v1951obus[temp_w*1 +:temp_w];
assign v1951ibus[data_w*1 +:data_w] = c799obus[data_w*5 +:data_w];
assign c799ibus[temp_w*6 +:temp_w] = v2047obus[temp_w*0 +:temp_w];
assign v2047ibus[data_w*0 +:data_w] = c799obus[data_w*6 +:data_w];
assign c800ibus[temp_w*0 +:temp_w] = v44obus[temp_w*1 +:temp_w];
assign v44ibus[data_w*1 +:data_w] = c800obus[data_w*0 +:data_w];
assign c800ibus[temp_w*1 +:temp_w] = v403obus[temp_w*2 +:temp_w];
assign v403ibus[data_w*2 +:data_w] = c800obus[data_w*1 +:data_w];
assign c800ibus[temp_w*2 +:temp_w] = v536obus[temp_w*3 +:temp_w];
assign v536ibus[data_w*3 +:data_w] = c800obus[data_w*2 +:data_w];
assign c800ibus[temp_w*3 +:temp_w] = v747obus[temp_w*3 +:temp_w];
assign v747ibus[data_w*3 +:data_w] = c800obus[data_w*3 +:data_w];
assign c800ibus[temp_w*4 +:temp_w] = v1139obus[temp_w*3 +:temp_w];
assign v1139ibus[data_w*3 +:data_w] = c800obus[data_w*4 +:data_w];
assign c800ibus[temp_w*5 +:temp_w] = v1952obus[temp_w*1 +:temp_w];
assign v1952ibus[data_w*1 +:data_w] = c800obus[data_w*5 +:data_w];
assign c800ibus[temp_w*6 +:temp_w] = v2048obus[temp_w*0 +:temp_w];
assign v2048ibus[data_w*0 +:data_w] = c800obus[data_w*6 +:data_w];
assign c801ibus[temp_w*0 +:temp_w] = v45obus[temp_w*1 +:temp_w];
assign v45ibus[data_w*1 +:data_w] = c801obus[data_w*0 +:data_w];
assign c801ibus[temp_w*1 +:temp_w] = v404obus[temp_w*2 +:temp_w];
assign v404ibus[data_w*2 +:data_w] = c801obus[data_w*1 +:data_w];
assign c801ibus[temp_w*2 +:temp_w] = v537obus[temp_w*3 +:temp_w];
assign v537ibus[data_w*3 +:data_w] = c801obus[data_w*2 +:data_w];
assign c801ibus[temp_w*3 +:temp_w] = v748obus[temp_w*3 +:temp_w];
assign v748ibus[data_w*3 +:data_w] = c801obus[data_w*3 +:data_w];
assign c801ibus[temp_w*4 +:temp_w] = v1140obus[temp_w*3 +:temp_w];
assign v1140ibus[data_w*3 +:data_w] = c801obus[data_w*4 +:data_w];
assign c801ibus[temp_w*5 +:temp_w] = v1953obus[temp_w*1 +:temp_w];
assign v1953ibus[data_w*1 +:data_w] = c801obus[data_w*5 +:data_w];
assign c801ibus[temp_w*6 +:temp_w] = v2049obus[temp_w*0 +:temp_w];
assign v2049ibus[data_w*0 +:data_w] = c801obus[data_w*6 +:data_w];
assign c802ibus[temp_w*0 +:temp_w] = v46obus[temp_w*1 +:temp_w];
assign v46ibus[data_w*1 +:data_w] = c802obus[data_w*0 +:data_w];
assign c802ibus[temp_w*1 +:temp_w] = v405obus[temp_w*2 +:temp_w];
assign v405ibus[data_w*2 +:data_w] = c802obus[data_w*1 +:data_w];
assign c802ibus[temp_w*2 +:temp_w] = v538obus[temp_w*3 +:temp_w];
assign v538ibus[data_w*3 +:data_w] = c802obus[data_w*2 +:data_w];
assign c802ibus[temp_w*3 +:temp_w] = v749obus[temp_w*3 +:temp_w];
assign v749ibus[data_w*3 +:data_w] = c802obus[data_w*3 +:data_w];
assign c802ibus[temp_w*4 +:temp_w] = v1141obus[temp_w*3 +:temp_w];
assign v1141ibus[data_w*3 +:data_w] = c802obus[data_w*4 +:data_w];
assign c802ibus[temp_w*5 +:temp_w] = v1954obus[temp_w*1 +:temp_w];
assign v1954ibus[data_w*1 +:data_w] = c802obus[data_w*5 +:data_w];
assign c802ibus[temp_w*6 +:temp_w] = v2050obus[temp_w*0 +:temp_w];
assign v2050ibus[data_w*0 +:data_w] = c802obus[data_w*6 +:data_w];
assign c803ibus[temp_w*0 +:temp_w] = v47obus[temp_w*1 +:temp_w];
assign v47ibus[data_w*1 +:data_w] = c803obus[data_w*0 +:data_w];
assign c803ibus[temp_w*1 +:temp_w] = v406obus[temp_w*2 +:temp_w];
assign v406ibus[data_w*2 +:data_w] = c803obus[data_w*1 +:data_w];
assign c803ibus[temp_w*2 +:temp_w] = v539obus[temp_w*3 +:temp_w];
assign v539ibus[data_w*3 +:data_w] = c803obus[data_w*2 +:data_w];
assign c803ibus[temp_w*3 +:temp_w] = v750obus[temp_w*3 +:temp_w];
assign v750ibus[data_w*3 +:data_w] = c803obus[data_w*3 +:data_w];
assign c803ibus[temp_w*4 +:temp_w] = v1142obus[temp_w*3 +:temp_w];
assign v1142ibus[data_w*3 +:data_w] = c803obus[data_w*4 +:data_w];
assign c803ibus[temp_w*5 +:temp_w] = v1955obus[temp_w*1 +:temp_w];
assign v1955ibus[data_w*1 +:data_w] = c803obus[data_w*5 +:data_w];
assign c803ibus[temp_w*6 +:temp_w] = v2051obus[temp_w*0 +:temp_w];
assign v2051ibus[data_w*0 +:data_w] = c803obus[data_w*6 +:data_w];
assign c804ibus[temp_w*0 +:temp_w] = v48obus[temp_w*1 +:temp_w];
assign v48ibus[data_w*1 +:data_w] = c804obus[data_w*0 +:data_w];
assign c804ibus[temp_w*1 +:temp_w] = v407obus[temp_w*2 +:temp_w];
assign v407ibus[data_w*2 +:data_w] = c804obus[data_w*1 +:data_w];
assign c804ibus[temp_w*2 +:temp_w] = v540obus[temp_w*3 +:temp_w];
assign v540ibus[data_w*3 +:data_w] = c804obus[data_w*2 +:data_w];
assign c804ibus[temp_w*3 +:temp_w] = v751obus[temp_w*3 +:temp_w];
assign v751ibus[data_w*3 +:data_w] = c804obus[data_w*3 +:data_w];
assign c804ibus[temp_w*4 +:temp_w] = v1143obus[temp_w*3 +:temp_w];
assign v1143ibus[data_w*3 +:data_w] = c804obus[data_w*4 +:data_w];
assign c804ibus[temp_w*5 +:temp_w] = v1956obus[temp_w*1 +:temp_w];
assign v1956ibus[data_w*1 +:data_w] = c804obus[data_w*5 +:data_w];
assign c804ibus[temp_w*6 +:temp_w] = v2052obus[temp_w*0 +:temp_w];
assign v2052ibus[data_w*0 +:data_w] = c804obus[data_w*6 +:data_w];
assign c805ibus[temp_w*0 +:temp_w] = v49obus[temp_w*1 +:temp_w];
assign v49ibus[data_w*1 +:data_w] = c805obus[data_w*0 +:data_w];
assign c805ibus[temp_w*1 +:temp_w] = v408obus[temp_w*2 +:temp_w];
assign v408ibus[data_w*2 +:data_w] = c805obus[data_w*1 +:data_w];
assign c805ibus[temp_w*2 +:temp_w] = v541obus[temp_w*3 +:temp_w];
assign v541ibus[data_w*3 +:data_w] = c805obus[data_w*2 +:data_w];
assign c805ibus[temp_w*3 +:temp_w] = v752obus[temp_w*3 +:temp_w];
assign v752ibus[data_w*3 +:data_w] = c805obus[data_w*3 +:data_w];
assign c805ibus[temp_w*4 +:temp_w] = v1144obus[temp_w*3 +:temp_w];
assign v1144ibus[data_w*3 +:data_w] = c805obus[data_w*4 +:data_w];
assign c805ibus[temp_w*5 +:temp_w] = v1957obus[temp_w*1 +:temp_w];
assign v1957ibus[data_w*1 +:data_w] = c805obus[data_w*5 +:data_w];
assign c805ibus[temp_w*6 +:temp_w] = v2053obus[temp_w*0 +:temp_w];
assign v2053ibus[data_w*0 +:data_w] = c805obus[data_w*6 +:data_w];
assign c806ibus[temp_w*0 +:temp_w] = v50obus[temp_w*1 +:temp_w];
assign v50ibus[data_w*1 +:data_w] = c806obus[data_w*0 +:data_w];
assign c806ibus[temp_w*1 +:temp_w] = v409obus[temp_w*2 +:temp_w];
assign v409ibus[data_w*2 +:data_w] = c806obus[data_w*1 +:data_w];
assign c806ibus[temp_w*2 +:temp_w] = v542obus[temp_w*3 +:temp_w];
assign v542ibus[data_w*3 +:data_w] = c806obus[data_w*2 +:data_w];
assign c806ibus[temp_w*3 +:temp_w] = v753obus[temp_w*3 +:temp_w];
assign v753ibus[data_w*3 +:data_w] = c806obus[data_w*3 +:data_w];
assign c806ibus[temp_w*4 +:temp_w] = v1145obus[temp_w*3 +:temp_w];
assign v1145ibus[data_w*3 +:data_w] = c806obus[data_w*4 +:data_w];
assign c806ibus[temp_w*5 +:temp_w] = v1958obus[temp_w*1 +:temp_w];
assign v1958ibus[data_w*1 +:data_w] = c806obus[data_w*5 +:data_w];
assign c806ibus[temp_w*6 +:temp_w] = v2054obus[temp_w*0 +:temp_w];
assign v2054ibus[data_w*0 +:data_w] = c806obus[data_w*6 +:data_w];
assign c807ibus[temp_w*0 +:temp_w] = v51obus[temp_w*1 +:temp_w];
assign v51ibus[data_w*1 +:data_w] = c807obus[data_w*0 +:data_w];
assign c807ibus[temp_w*1 +:temp_w] = v410obus[temp_w*2 +:temp_w];
assign v410ibus[data_w*2 +:data_w] = c807obus[data_w*1 +:data_w];
assign c807ibus[temp_w*2 +:temp_w] = v543obus[temp_w*3 +:temp_w];
assign v543ibus[data_w*3 +:data_w] = c807obus[data_w*2 +:data_w];
assign c807ibus[temp_w*3 +:temp_w] = v754obus[temp_w*3 +:temp_w];
assign v754ibus[data_w*3 +:data_w] = c807obus[data_w*3 +:data_w];
assign c807ibus[temp_w*4 +:temp_w] = v1146obus[temp_w*3 +:temp_w];
assign v1146ibus[data_w*3 +:data_w] = c807obus[data_w*4 +:data_w];
assign c807ibus[temp_w*5 +:temp_w] = v1959obus[temp_w*1 +:temp_w];
assign v1959ibus[data_w*1 +:data_w] = c807obus[data_w*5 +:data_w];
assign c807ibus[temp_w*6 +:temp_w] = v2055obus[temp_w*0 +:temp_w];
assign v2055ibus[data_w*0 +:data_w] = c807obus[data_w*6 +:data_w];
assign c808ibus[temp_w*0 +:temp_w] = v52obus[temp_w*1 +:temp_w];
assign v52ibus[data_w*1 +:data_w] = c808obus[data_w*0 +:data_w];
assign c808ibus[temp_w*1 +:temp_w] = v411obus[temp_w*2 +:temp_w];
assign v411ibus[data_w*2 +:data_w] = c808obus[data_w*1 +:data_w];
assign c808ibus[temp_w*2 +:temp_w] = v544obus[temp_w*3 +:temp_w];
assign v544ibus[data_w*3 +:data_w] = c808obus[data_w*2 +:data_w];
assign c808ibus[temp_w*3 +:temp_w] = v755obus[temp_w*3 +:temp_w];
assign v755ibus[data_w*3 +:data_w] = c808obus[data_w*3 +:data_w];
assign c808ibus[temp_w*4 +:temp_w] = v1147obus[temp_w*3 +:temp_w];
assign v1147ibus[data_w*3 +:data_w] = c808obus[data_w*4 +:data_w];
assign c808ibus[temp_w*5 +:temp_w] = v1960obus[temp_w*1 +:temp_w];
assign v1960ibus[data_w*1 +:data_w] = c808obus[data_w*5 +:data_w];
assign c808ibus[temp_w*6 +:temp_w] = v2056obus[temp_w*0 +:temp_w];
assign v2056ibus[data_w*0 +:data_w] = c808obus[data_w*6 +:data_w];
assign c809ibus[temp_w*0 +:temp_w] = v53obus[temp_w*1 +:temp_w];
assign v53ibus[data_w*1 +:data_w] = c809obus[data_w*0 +:data_w];
assign c809ibus[temp_w*1 +:temp_w] = v412obus[temp_w*2 +:temp_w];
assign v412ibus[data_w*2 +:data_w] = c809obus[data_w*1 +:data_w];
assign c809ibus[temp_w*2 +:temp_w] = v545obus[temp_w*3 +:temp_w];
assign v545ibus[data_w*3 +:data_w] = c809obus[data_w*2 +:data_w];
assign c809ibus[temp_w*3 +:temp_w] = v756obus[temp_w*3 +:temp_w];
assign v756ibus[data_w*3 +:data_w] = c809obus[data_w*3 +:data_w];
assign c809ibus[temp_w*4 +:temp_w] = v1148obus[temp_w*3 +:temp_w];
assign v1148ibus[data_w*3 +:data_w] = c809obus[data_w*4 +:data_w];
assign c809ibus[temp_w*5 +:temp_w] = v1961obus[temp_w*1 +:temp_w];
assign v1961ibus[data_w*1 +:data_w] = c809obus[data_w*5 +:data_w];
assign c809ibus[temp_w*6 +:temp_w] = v2057obus[temp_w*0 +:temp_w];
assign v2057ibus[data_w*0 +:data_w] = c809obus[data_w*6 +:data_w];
assign c810ibus[temp_w*0 +:temp_w] = v54obus[temp_w*1 +:temp_w];
assign v54ibus[data_w*1 +:data_w] = c810obus[data_w*0 +:data_w];
assign c810ibus[temp_w*1 +:temp_w] = v413obus[temp_w*2 +:temp_w];
assign v413ibus[data_w*2 +:data_w] = c810obus[data_w*1 +:data_w];
assign c810ibus[temp_w*2 +:temp_w] = v546obus[temp_w*3 +:temp_w];
assign v546ibus[data_w*3 +:data_w] = c810obus[data_w*2 +:data_w];
assign c810ibus[temp_w*3 +:temp_w] = v757obus[temp_w*3 +:temp_w];
assign v757ibus[data_w*3 +:data_w] = c810obus[data_w*3 +:data_w];
assign c810ibus[temp_w*4 +:temp_w] = v1149obus[temp_w*3 +:temp_w];
assign v1149ibus[data_w*3 +:data_w] = c810obus[data_w*4 +:data_w];
assign c810ibus[temp_w*5 +:temp_w] = v1962obus[temp_w*1 +:temp_w];
assign v1962ibus[data_w*1 +:data_w] = c810obus[data_w*5 +:data_w];
assign c810ibus[temp_w*6 +:temp_w] = v2058obus[temp_w*0 +:temp_w];
assign v2058ibus[data_w*0 +:data_w] = c810obus[data_w*6 +:data_w];
assign c811ibus[temp_w*0 +:temp_w] = v55obus[temp_w*1 +:temp_w];
assign v55ibus[data_w*1 +:data_w] = c811obus[data_w*0 +:data_w];
assign c811ibus[temp_w*1 +:temp_w] = v414obus[temp_w*2 +:temp_w];
assign v414ibus[data_w*2 +:data_w] = c811obus[data_w*1 +:data_w];
assign c811ibus[temp_w*2 +:temp_w] = v547obus[temp_w*3 +:temp_w];
assign v547ibus[data_w*3 +:data_w] = c811obus[data_w*2 +:data_w];
assign c811ibus[temp_w*3 +:temp_w] = v758obus[temp_w*3 +:temp_w];
assign v758ibus[data_w*3 +:data_w] = c811obus[data_w*3 +:data_w];
assign c811ibus[temp_w*4 +:temp_w] = v1150obus[temp_w*3 +:temp_w];
assign v1150ibus[data_w*3 +:data_w] = c811obus[data_w*4 +:data_w];
assign c811ibus[temp_w*5 +:temp_w] = v1963obus[temp_w*1 +:temp_w];
assign v1963ibus[data_w*1 +:data_w] = c811obus[data_w*5 +:data_w];
assign c811ibus[temp_w*6 +:temp_w] = v2059obus[temp_w*0 +:temp_w];
assign v2059ibus[data_w*0 +:data_w] = c811obus[data_w*6 +:data_w];
assign c812ibus[temp_w*0 +:temp_w] = v56obus[temp_w*1 +:temp_w];
assign v56ibus[data_w*1 +:data_w] = c812obus[data_w*0 +:data_w];
assign c812ibus[temp_w*1 +:temp_w] = v415obus[temp_w*2 +:temp_w];
assign v415ibus[data_w*2 +:data_w] = c812obus[data_w*1 +:data_w];
assign c812ibus[temp_w*2 +:temp_w] = v548obus[temp_w*3 +:temp_w];
assign v548ibus[data_w*3 +:data_w] = c812obus[data_w*2 +:data_w];
assign c812ibus[temp_w*3 +:temp_w] = v759obus[temp_w*3 +:temp_w];
assign v759ibus[data_w*3 +:data_w] = c812obus[data_w*3 +:data_w];
assign c812ibus[temp_w*4 +:temp_w] = v1151obus[temp_w*3 +:temp_w];
assign v1151ibus[data_w*3 +:data_w] = c812obus[data_w*4 +:data_w];
assign c812ibus[temp_w*5 +:temp_w] = v1964obus[temp_w*1 +:temp_w];
assign v1964ibus[data_w*1 +:data_w] = c812obus[data_w*5 +:data_w];
assign c812ibus[temp_w*6 +:temp_w] = v2060obus[temp_w*0 +:temp_w];
assign v2060ibus[data_w*0 +:data_w] = c812obus[data_w*6 +:data_w];
assign c813ibus[temp_w*0 +:temp_w] = v57obus[temp_w*1 +:temp_w];
assign v57ibus[data_w*1 +:data_w] = c813obus[data_w*0 +:data_w];
assign c813ibus[temp_w*1 +:temp_w] = v416obus[temp_w*2 +:temp_w];
assign v416ibus[data_w*2 +:data_w] = c813obus[data_w*1 +:data_w];
assign c813ibus[temp_w*2 +:temp_w] = v549obus[temp_w*3 +:temp_w];
assign v549ibus[data_w*3 +:data_w] = c813obus[data_w*2 +:data_w];
assign c813ibus[temp_w*3 +:temp_w] = v760obus[temp_w*3 +:temp_w];
assign v760ibus[data_w*3 +:data_w] = c813obus[data_w*3 +:data_w];
assign c813ibus[temp_w*4 +:temp_w] = v1056obus[temp_w*3 +:temp_w];
assign v1056ibus[data_w*3 +:data_w] = c813obus[data_w*4 +:data_w];
assign c813ibus[temp_w*5 +:temp_w] = v1965obus[temp_w*1 +:temp_w];
assign v1965ibus[data_w*1 +:data_w] = c813obus[data_w*5 +:data_w];
assign c813ibus[temp_w*6 +:temp_w] = v2061obus[temp_w*0 +:temp_w];
assign v2061ibus[data_w*0 +:data_w] = c813obus[data_w*6 +:data_w];
assign c814ibus[temp_w*0 +:temp_w] = v58obus[temp_w*1 +:temp_w];
assign v58ibus[data_w*1 +:data_w] = c814obus[data_w*0 +:data_w];
assign c814ibus[temp_w*1 +:temp_w] = v417obus[temp_w*2 +:temp_w];
assign v417ibus[data_w*2 +:data_w] = c814obus[data_w*1 +:data_w];
assign c814ibus[temp_w*2 +:temp_w] = v550obus[temp_w*3 +:temp_w];
assign v550ibus[data_w*3 +:data_w] = c814obus[data_w*2 +:data_w];
assign c814ibus[temp_w*3 +:temp_w] = v761obus[temp_w*3 +:temp_w];
assign v761ibus[data_w*3 +:data_w] = c814obus[data_w*3 +:data_w];
assign c814ibus[temp_w*4 +:temp_w] = v1057obus[temp_w*3 +:temp_w];
assign v1057ibus[data_w*3 +:data_w] = c814obus[data_w*4 +:data_w];
assign c814ibus[temp_w*5 +:temp_w] = v1966obus[temp_w*1 +:temp_w];
assign v1966ibus[data_w*1 +:data_w] = c814obus[data_w*5 +:data_w];
assign c814ibus[temp_w*6 +:temp_w] = v2062obus[temp_w*0 +:temp_w];
assign v2062ibus[data_w*0 +:data_w] = c814obus[data_w*6 +:data_w];
assign c815ibus[temp_w*0 +:temp_w] = v59obus[temp_w*1 +:temp_w];
assign v59ibus[data_w*1 +:data_w] = c815obus[data_w*0 +:data_w];
assign c815ibus[temp_w*1 +:temp_w] = v418obus[temp_w*2 +:temp_w];
assign v418ibus[data_w*2 +:data_w] = c815obus[data_w*1 +:data_w];
assign c815ibus[temp_w*2 +:temp_w] = v551obus[temp_w*3 +:temp_w];
assign v551ibus[data_w*3 +:data_w] = c815obus[data_w*2 +:data_w];
assign c815ibus[temp_w*3 +:temp_w] = v762obus[temp_w*3 +:temp_w];
assign v762ibus[data_w*3 +:data_w] = c815obus[data_w*3 +:data_w];
assign c815ibus[temp_w*4 +:temp_w] = v1058obus[temp_w*3 +:temp_w];
assign v1058ibus[data_w*3 +:data_w] = c815obus[data_w*4 +:data_w];
assign c815ibus[temp_w*5 +:temp_w] = v1967obus[temp_w*1 +:temp_w];
assign v1967ibus[data_w*1 +:data_w] = c815obus[data_w*5 +:data_w];
assign c815ibus[temp_w*6 +:temp_w] = v2063obus[temp_w*0 +:temp_w];
assign v2063ibus[data_w*0 +:data_w] = c815obus[data_w*6 +:data_w];
assign c816ibus[temp_w*0 +:temp_w] = v60obus[temp_w*1 +:temp_w];
assign v60ibus[data_w*1 +:data_w] = c816obus[data_w*0 +:data_w];
assign c816ibus[temp_w*1 +:temp_w] = v419obus[temp_w*2 +:temp_w];
assign v419ibus[data_w*2 +:data_w] = c816obus[data_w*1 +:data_w];
assign c816ibus[temp_w*2 +:temp_w] = v552obus[temp_w*3 +:temp_w];
assign v552ibus[data_w*3 +:data_w] = c816obus[data_w*2 +:data_w];
assign c816ibus[temp_w*3 +:temp_w] = v763obus[temp_w*3 +:temp_w];
assign v763ibus[data_w*3 +:data_w] = c816obus[data_w*3 +:data_w];
assign c816ibus[temp_w*4 +:temp_w] = v1059obus[temp_w*3 +:temp_w];
assign v1059ibus[data_w*3 +:data_w] = c816obus[data_w*4 +:data_w];
assign c816ibus[temp_w*5 +:temp_w] = v1968obus[temp_w*1 +:temp_w];
assign v1968ibus[data_w*1 +:data_w] = c816obus[data_w*5 +:data_w];
assign c816ibus[temp_w*6 +:temp_w] = v2064obus[temp_w*0 +:temp_w];
assign v2064ibus[data_w*0 +:data_w] = c816obus[data_w*6 +:data_w];
assign c817ibus[temp_w*0 +:temp_w] = v61obus[temp_w*1 +:temp_w];
assign v61ibus[data_w*1 +:data_w] = c817obus[data_w*0 +:data_w];
assign c817ibus[temp_w*1 +:temp_w] = v420obus[temp_w*2 +:temp_w];
assign v420ibus[data_w*2 +:data_w] = c817obus[data_w*1 +:data_w];
assign c817ibus[temp_w*2 +:temp_w] = v553obus[temp_w*3 +:temp_w];
assign v553ibus[data_w*3 +:data_w] = c817obus[data_w*2 +:data_w];
assign c817ibus[temp_w*3 +:temp_w] = v764obus[temp_w*3 +:temp_w];
assign v764ibus[data_w*3 +:data_w] = c817obus[data_w*3 +:data_w];
assign c817ibus[temp_w*4 +:temp_w] = v1060obus[temp_w*3 +:temp_w];
assign v1060ibus[data_w*3 +:data_w] = c817obus[data_w*4 +:data_w];
assign c817ibus[temp_w*5 +:temp_w] = v1969obus[temp_w*1 +:temp_w];
assign v1969ibus[data_w*1 +:data_w] = c817obus[data_w*5 +:data_w];
assign c817ibus[temp_w*6 +:temp_w] = v2065obus[temp_w*0 +:temp_w];
assign v2065ibus[data_w*0 +:data_w] = c817obus[data_w*6 +:data_w];
assign c818ibus[temp_w*0 +:temp_w] = v62obus[temp_w*1 +:temp_w];
assign v62ibus[data_w*1 +:data_w] = c818obus[data_w*0 +:data_w];
assign c818ibus[temp_w*1 +:temp_w] = v421obus[temp_w*2 +:temp_w];
assign v421ibus[data_w*2 +:data_w] = c818obus[data_w*1 +:data_w];
assign c818ibus[temp_w*2 +:temp_w] = v554obus[temp_w*3 +:temp_w];
assign v554ibus[data_w*3 +:data_w] = c818obus[data_w*2 +:data_w];
assign c818ibus[temp_w*3 +:temp_w] = v765obus[temp_w*3 +:temp_w];
assign v765ibus[data_w*3 +:data_w] = c818obus[data_w*3 +:data_w];
assign c818ibus[temp_w*4 +:temp_w] = v1061obus[temp_w*3 +:temp_w];
assign v1061ibus[data_w*3 +:data_w] = c818obus[data_w*4 +:data_w];
assign c818ibus[temp_w*5 +:temp_w] = v1970obus[temp_w*1 +:temp_w];
assign v1970ibus[data_w*1 +:data_w] = c818obus[data_w*5 +:data_w];
assign c818ibus[temp_w*6 +:temp_w] = v2066obus[temp_w*0 +:temp_w];
assign v2066ibus[data_w*0 +:data_w] = c818obus[data_w*6 +:data_w];
assign c819ibus[temp_w*0 +:temp_w] = v63obus[temp_w*1 +:temp_w];
assign v63ibus[data_w*1 +:data_w] = c819obus[data_w*0 +:data_w];
assign c819ibus[temp_w*1 +:temp_w] = v422obus[temp_w*2 +:temp_w];
assign v422ibus[data_w*2 +:data_w] = c819obus[data_w*1 +:data_w];
assign c819ibus[temp_w*2 +:temp_w] = v555obus[temp_w*3 +:temp_w];
assign v555ibus[data_w*3 +:data_w] = c819obus[data_w*2 +:data_w];
assign c819ibus[temp_w*3 +:temp_w] = v766obus[temp_w*3 +:temp_w];
assign v766ibus[data_w*3 +:data_w] = c819obus[data_w*3 +:data_w];
assign c819ibus[temp_w*4 +:temp_w] = v1062obus[temp_w*3 +:temp_w];
assign v1062ibus[data_w*3 +:data_w] = c819obus[data_w*4 +:data_w];
assign c819ibus[temp_w*5 +:temp_w] = v1971obus[temp_w*1 +:temp_w];
assign v1971ibus[data_w*1 +:data_w] = c819obus[data_w*5 +:data_w];
assign c819ibus[temp_w*6 +:temp_w] = v2067obus[temp_w*0 +:temp_w];
assign v2067ibus[data_w*0 +:data_w] = c819obus[data_w*6 +:data_w];
assign c820ibus[temp_w*0 +:temp_w] = v64obus[temp_w*1 +:temp_w];
assign v64ibus[data_w*1 +:data_w] = c820obus[data_w*0 +:data_w];
assign c820ibus[temp_w*1 +:temp_w] = v423obus[temp_w*2 +:temp_w];
assign v423ibus[data_w*2 +:data_w] = c820obus[data_w*1 +:data_w];
assign c820ibus[temp_w*2 +:temp_w] = v556obus[temp_w*3 +:temp_w];
assign v556ibus[data_w*3 +:data_w] = c820obus[data_w*2 +:data_w];
assign c820ibus[temp_w*3 +:temp_w] = v767obus[temp_w*3 +:temp_w];
assign v767ibus[data_w*3 +:data_w] = c820obus[data_w*3 +:data_w];
assign c820ibus[temp_w*4 +:temp_w] = v1063obus[temp_w*3 +:temp_w];
assign v1063ibus[data_w*3 +:data_w] = c820obus[data_w*4 +:data_w];
assign c820ibus[temp_w*5 +:temp_w] = v1972obus[temp_w*1 +:temp_w];
assign v1972ibus[data_w*1 +:data_w] = c820obus[data_w*5 +:data_w];
assign c820ibus[temp_w*6 +:temp_w] = v2068obus[temp_w*0 +:temp_w];
assign v2068ibus[data_w*0 +:data_w] = c820obus[data_w*6 +:data_w];
assign c821ibus[temp_w*0 +:temp_w] = v65obus[temp_w*1 +:temp_w];
assign v65ibus[data_w*1 +:data_w] = c821obus[data_w*0 +:data_w];
assign c821ibus[temp_w*1 +:temp_w] = v424obus[temp_w*2 +:temp_w];
assign v424ibus[data_w*2 +:data_w] = c821obus[data_w*1 +:data_w];
assign c821ibus[temp_w*2 +:temp_w] = v557obus[temp_w*3 +:temp_w];
assign v557ibus[data_w*3 +:data_w] = c821obus[data_w*2 +:data_w];
assign c821ibus[temp_w*3 +:temp_w] = v672obus[temp_w*3 +:temp_w];
assign v672ibus[data_w*3 +:data_w] = c821obus[data_w*3 +:data_w];
assign c821ibus[temp_w*4 +:temp_w] = v1064obus[temp_w*3 +:temp_w];
assign v1064ibus[data_w*3 +:data_w] = c821obus[data_w*4 +:data_w];
assign c821ibus[temp_w*5 +:temp_w] = v1973obus[temp_w*1 +:temp_w];
assign v1973ibus[data_w*1 +:data_w] = c821obus[data_w*5 +:data_w];
assign c821ibus[temp_w*6 +:temp_w] = v2069obus[temp_w*0 +:temp_w];
assign v2069ibus[data_w*0 +:data_w] = c821obus[data_w*6 +:data_w];
assign c822ibus[temp_w*0 +:temp_w] = v66obus[temp_w*1 +:temp_w];
assign v66ibus[data_w*1 +:data_w] = c822obus[data_w*0 +:data_w];
assign c822ibus[temp_w*1 +:temp_w] = v425obus[temp_w*2 +:temp_w];
assign v425ibus[data_w*2 +:data_w] = c822obus[data_w*1 +:data_w];
assign c822ibus[temp_w*2 +:temp_w] = v558obus[temp_w*3 +:temp_w];
assign v558ibus[data_w*3 +:data_w] = c822obus[data_w*2 +:data_w];
assign c822ibus[temp_w*3 +:temp_w] = v673obus[temp_w*3 +:temp_w];
assign v673ibus[data_w*3 +:data_w] = c822obus[data_w*3 +:data_w];
assign c822ibus[temp_w*4 +:temp_w] = v1065obus[temp_w*3 +:temp_w];
assign v1065ibus[data_w*3 +:data_w] = c822obus[data_w*4 +:data_w];
assign c822ibus[temp_w*5 +:temp_w] = v1974obus[temp_w*1 +:temp_w];
assign v1974ibus[data_w*1 +:data_w] = c822obus[data_w*5 +:data_w];
assign c822ibus[temp_w*6 +:temp_w] = v2070obus[temp_w*0 +:temp_w];
assign v2070ibus[data_w*0 +:data_w] = c822obus[data_w*6 +:data_w];
assign c823ibus[temp_w*0 +:temp_w] = v67obus[temp_w*1 +:temp_w];
assign v67ibus[data_w*1 +:data_w] = c823obus[data_w*0 +:data_w];
assign c823ibus[temp_w*1 +:temp_w] = v426obus[temp_w*2 +:temp_w];
assign v426ibus[data_w*2 +:data_w] = c823obus[data_w*1 +:data_w];
assign c823ibus[temp_w*2 +:temp_w] = v559obus[temp_w*3 +:temp_w];
assign v559ibus[data_w*3 +:data_w] = c823obus[data_w*2 +:data_w];
assign c823ibus[temp_w*3 +:temp_w] = v674obus[temp_w*3 +:temp_w];
assign v674ibus[data_w*3 +:data_w] = c823obus[data_w*3 +:data_w];
assign c823ibus[temp_w*4 +:temp_w] = v1066obus[temp_w*3 +:temp_w];
assign v1066ibus[data_w*3 +:data_w] = c823obus[data_w*4 +:data_w];
assign c823ibus[temp_w*5 +:temp_w] = v1975obus[temp_w*1 +:temp_w];
assign v1975ibus[data_w*1 +:data_w] = c823obus[data_w*5 +:data_w];
assign c823ibus[temp_w*6 +:temp_w] = v2071obus[temp_w*0 +:temp_w];
assign v2071ibus[data_w*0 +:data_w] = c823obus[data_w*6 +:data_w];
assign c824ibus[temp_w*0 +:temp_w] = v68obus[temp_w*1 +:temp_w];
assign v68ibus[data_w*1 +:data_w] = c824obus[data_w*0 +:data_w];
assign c824ibus[temp_w*1 +:temp_w] = v427obus[temp_w*2 +:temp_w];
assign v427ibus[data_w*2 +:data_w] = c824obus[data_w*1 +:data_w];
assign c824ibus[temp_w*2 +:temp_w] = v560obus[temp_w*3 +:temp_w];
assign v560ibus[data_w*3 +:data_w] = c824obus[data_w*2 +:data_w];
assign c824ibus[temp_w*3 +:temp_w] = v675obus[temp_w*3 +:temp_w];
assign v675ibus[data_w*3 +:data_w] = c824obus[data_w*3 +:data_w];
assign c824ibus[temp_w*4 +:temp_w] = v1067obus[temp_w*3 +:temp_w];
assign v1067ibus[data_w*3 +:data_w] = c824obus[data_w*4 +:data_w];
assign c824ibus[temp_w*5 +:temp_w] = v1976obus[temp_w*1 +:temp_w];
assign v1976ibus[data_w*1 +:data_w] = c824obus[data_w*5 +:data_w];
assign c824ibus[temp_w*6 +:temp_w] = v2072obus[temp_w*0 +:temp_w];
assign v2072ibus[data_w*0 +:data_w] = c824obus[data_w*6 +:data_w];
assign c825ibus[temp_w*0 +:temp_w] = v69obus[temp_w*1 +:temp_w];
assign v69ibus[data_w*1 +:data_w] = c825obus[data_w*0 +:data_w];
assign c825ibus[temp_w*1 +:temp_w] = v428obus[temp_w*2 +:temp_w];
assign v428ibus[data_w*2 +:data_w] = c825obus[data_w*1 +:data_w];
assign c825ibus[temp_w*2 +:temp_w] = v561obus[temp_w*3 +:temp_w];
assign v561ibus[data_w*3 +:data_w] = c825obus[data_w*2 +:data_w];
assign c825ibus[temp_w*3 +:temp_w] = v676obus[temp_w*3 +:temp_w];
assign v676ibus[data_w*3 +:data_w] = c825obus[data_w*3 +:data_w];
assign c825ibus[temp_w*4 +:temp_w] = v1068obus[temp_w*3 +:temp_w];
assign v1068ibus[data_w*3 +:data_w] = c825obus[data_w*4 +:data_w];
assign c825ibus[temp_w*5 +:temp_w] = v1977obus[temp_w*1 +:temp_w];
assign v1977ibus[data_w*1 +:data_w] = c825obus[data_w*5 +:data_w];
assign c825ibus[temp_w*6 +:temp_w] = v2073obus[temp_w*0 +:temp_w];
assign v2073ibus[data_w*0 +:data_w] = c825obus[data_w*6 +:data_w];
assign c826ibus[temp_w*0 +:temp_w] = v70obus[temp_w*1 +:temp_w];
assign v70ibus[data_w*1 +:data_w] = c826obus[data_w*0 +:data_w];
assign c826ibus[temp_w*1 +:temp_w] = v429obus[temp_w*2 +:temp_w];
assign v429ibus[data_w*2 +:data_w] = c826obus[data_w*1 +:data_w];
assign c826ibus[temp_w*2 +:temp_w] = v562obus[temp_w*3 +:temp_w];
assign v562ibus[data_w*3 +:data_w] = c826obus[data_w*2 +:data_w];
assign c826ibus[temp_w*3 +:temp_w] = v677obus[temp_w*3 +:temp_w];
assign v677ibus[data_w*3 +:data_w] = c826obus[data_w*3 +:data_w];
assign c826ibus[temp_w*4 +:temp_w] = v1069obus[temp_w*3 +:temp_w];
assign v1069ibus[data_w*3 +:data_w] = c826obus[data_w*4 +:data_w];
assign c826ibus[temp_w*5 +:temp_w] = v1978obus[temp_w*1 +:temp_w];
assign v1978ibus[data_w*1 +:data_w] = c826obus[data_w*5 +:data_w];
assign c826ibus[temp_w*6 +:temp_w] = v2074obus[temp_w*0 +:temp_w];
assign v2074ibus[data_w*0 +:data_w] = c826obus[data_w*6 +:data_w];
assign c827ibus[temp_w*0 +:temp_w] = v71obus[temp_w*1 +:temp_w];
assign v71ibus[data_w*1 +:data_w] = c827obus[data_w*0 +:data_w];
assign c827ibus[temp_w*1 +:temp_w] = v430obus[temp_w*2 +:temp_w];
assign v430ibus[data_w*2 +:data_w] = c827obus[data_w*1 +:data_w];
assign c827ibus[temp_w*2 +:temp_w] = v563obus[temp_w*3 +:temp_w];
assign v563ibus[data_w*3 +:data_w] = c827obus[data_w*2 +:data_w];
assign c827ibus[temp_w*3 +:temp_w] = v678obus[temp_w*3 +:temp_w];
assign v678ibus[data_w*3 +:data_w] = c827obus[data_w*3 +:data_w];
assign c827ibus[temp_w*4 +:temp_w] = v1070obus[temp_w*3 +:temp_w];
assign v1070ibus[data_w*3 +:data_w] = c827obus[data_w*4 +:data_w];
assign c827ibus[temp_w*5 +:temp_w] = v1979obus[temp_w*1 +:temp_w];
assign v1979ibus[data_w*1 +:data_w] = c827obus[data_w*5 +:data_w];
assign c827ibus[temp_w*6 +:temp_w] = v2075obus[temp_w*0 +:temp_w];
assign v2075ibus[data_w*0 +:data_w] = c827obus[data_w*6 +:data_w];
assign c828ibus[temp_w*0 +:temp_w] = v72obus[temp_w*1 +:temp_w];
assign v72ibus[data_w*1 +:data_w] = c828obus[data_w*0 +:data_w];
assign c828ibus[temp_w*1 +:temp_w] = v431obus[temp_w*2 +:temp_w];
assign v431ibus[data_w*2 +:data_w] = c828obus[data_w*1 +:data_w];
assign c828ibus[temp_w*2 +:temp_w] = v564obus[temp_w*3 +:temp_w];
assign v564ibus[data_w*3 +:data_w] = c828obus[data_w*2 +:data_w];
assign c828ibus[temp_w*3 +:temp_w] = v679obus[temp_w*3 +:temp_w];
assign v679ibus[data_w*3 +:data_w] = c828obus[data_w*3 +:data_w];
assign c828ibus[temp_w*4 +:temp_w] = v1071obus[temp_w*3 +:temp_w];
assign v1071ibus[data_w*3 +:data_w] = c828obus[data_w*4 +:data_w];
assign c828ibus[temp_w*5 +:temp_w] = v1980obus[temp_w*1 +:temp_w];
assign v1980ibus[data_w*1 +:data_w] = c828obus[data_w*5 +:data_w];
assign c828ibus[temp_w*6 +:temp_w] = v2076obus[temp_w*0 +:temp_w];
assign v2076ibus[data_w*0 +:data_w] = c828obus[data_w*6 +:data_w];
assign c829ibus[temp_w*0 +:temp_w] = v73obus[temp_w*1 +:temp_w];
assign v73ibus[data_w*1 +:data_w] = c829obus[data_w*0 +:data_w];
assign c829ibus[temp_w*1 +:temp_w] = v432obus[temp_w*2 +:temp_w];
assign v432ibus[data_w*2 +:data_w] = c829obus[data_w*1 +:data_w];
assign c829ibus[temp_w*2 +:temp_w] = v565obus[temp_w*3 +:temp_w];
assign v565ibus[data_w*3 +:data_w] = c829obus[data_w*2 +:data_w];
assign c829ibus[temp_w*3 +:temp_w] = v680obus[temp_w*3 +:temp_w];
assign v680ibus[data_w*3 +:data_w] = c829obus[data_w*3 +:data_w];
assign c829ibus[temp_w*4 +:temp_w] = v1072obus[temp_w*3 +:temp_w];
assign v1072ibus[data_w*3 +:data_w] = c829obus[data_w*4 +:data_w];
assign c829ibus[temp_w*5 +:temp_w] = v1981obus[temp_w*1 +:temp_w];
assign v1981ibus[data_w*1 +:data_w] = c829obus[data_w*5 +:data_w];
assign c829ibus[temp_w*6 +:temp_w] = v2077obus[temp_w*0 +:temp_w];
assign v2077ibus[data_w*0 +:data_w] = c829obus[data_w*6 +:data_w];
assign c830ibus[temp_w*0 +:temp_w] = v74obus[temp_w*1 +:temp_w];
assign v74ibus[data_w*1 +:data_w] = c830obus[data_w*0 +:data_w];
assign c830ibus[temp_w*1 +:temp_w] = v433obus[temp_w*2 +:temp_w];
assign v433ibus[data_w*2 +:data_w] = c830obus[data_w*1 +:data_w];
assign c830ibus[temp_w*2 +:temp_w] = v566obus[temp_w*3 +:temp_w];
assign v566ibus[data_w*3 +:data_w] = c830obus[data_w*2 +:data_w];
assign c830ibus[temp_w*3 +:temp_w] = v681obus[temp_w*3 +:temp_w];
assign v681ibus[data_w*3 +:data_w] = c830obus[data_w*3 +:data_w];
assign c830ibus[temp_w*4 +:temp_w] = v1073obus[temp_w*3 +:temp_w];
assign v1073ibus[data_w*3 +:data_w] = c830obus[data_w*4 +:data_w];
assign c830ibus[temp_w*5 +:temp_w] = v1982obus[temp_w*1 +:temp_w];
assign v1982ibus[data_w*1 +:data_w] = c830obus[data_w*5 +:data_w];
assign c830ibus[temp_w*6 +:temp_w] = v2078obus[temp_w*0 +:temp_w];
assign v2078ibus[data_w*0 +:data_w] = c830obus[data_w*6 +:data_w];
assign c831ibus[temp_w*0 +:temp_w] = v75obus[temp_w*1 +:temp_w];
assign v75ibus[data_w*1 +:data_w] = c831obus[data_w*0 +:data_w];
assign c831ibus[temp_w*1 +:temp_w] = v434obus[temp_w*2 +:temp_w];
assign v434ibus[data_w*2 +:data_w] = c831obus[data_w*1 +:data_w];
assign c831ibus[temp_w*2 +:temp_w] = v567obus[temp_w*3 +:temp_w];
assign v567ibus[data_w*3 +:data_w] = c831obus[data_w*2 +:data_w];
assign c831ibus[temp_w*3 +:temp_w] = v682obus[temp_w*3 +:temp_w];
assign v682ibus[data_w*3 +:data_w] = c831obus[data_w*3 +:data_w];
assign c831ibus[temp_w*4 +:temp_w] = v1074obus[temp_w*3 +:temp_w];
assign v1074ibus[data_w*3 +:data_w] = c831obus[data_w*4 +:data_w];
assign c831ibus[temp_w*5 +:temp_w] = v1983obus[temp_w*1 +:temp_w];
assign v1983ibus[data_w*1 +:data_w] = c831obus[data_w*5 +:data_w];
assign c831ibus[temp_w*6 +:temp_w] = v2079obus[temp_w*0 +:temp_w];
assign v2079ibus[data_w*0 +:data_w] = c831obus[data_w*6 +:data_w];
assign c832ibus[temp_w*0 +:temp_w] = v76obus[temp_w*1 +:temp_w];
assign v76ibus[data_w*1 +:data_w] = c832obus[data_w*0 +:data_w];
assign c832ibus[temp_w*1 +:temp_w] = v435obus[temp_w*2 +:temp_w];
assign v435ibus[data_w*2 +:data_w] = c832obus[data_w*1 +:data_w];
assign c832ibus[temp_w*2 +:temp_w] = v568obus[temp_w*3 +:temp_w];
assign v568ibus[data_w*3 +:data_w] = c832obus[data_w*2 +:data_w];
assign c832ibus[temp_w*3 +:temp_w] = v683obus[temp_w*3 +:temp_w];
assign v683ibus[data_w*3 +:data_w] = c832obus[data_w*3 +:data_w];
assign c832ibus[temp_w*4 +:temp_w] = v1075obus[temp_w*3 +:temp_w];
assign v1075ibus[data_w*3 +:data_w] = c832obus[data_w*4 +:data_w];
assign c832ibus[temp_w*5 +:temp_w] = v1984obus[temp_w*1 +:temp_w];
assign v1984ibus[data_w*1 +:data_w] = c832obus[data_w*5 +:data_w];
assign c832ibus[temp_w*6 +:temp_w] = v2080obus[temp_w*0 +:temp_w];
assign v2080ibus[data_w*0 +:data_w] = c832obus[data_w*6 +:data_w];
assign c833ibus[temp_w*0 +:temp_w] = v77obus[temp_w*1 +:temp_w];
assign v77ibus[data_w*1 +:data_w] = c833obus[data_w*0 +:data_w];
assign c833ibus[temp_w*1 +:temp_w] = v436obus[temp_w*2 +:temp_w];
assign v436ibus[data_w*2 +:data_w] = c833obus[data_w*1 +:data_w];
assign c833ibus[temp_w*2 +:temp_w] = v569obus[temp_w*3 +:temp_w];
assign v569ibus[data_w*3 +:data_w] = c833obus[data_w*2 +:data_w];
assign c833ibus[temp_w*3 +:temp_w] = v684obus[temp_w*3 +:temp_w];
assign v684ibus[data_w*3 +:data_w] = c833obus[data_w*3 +:data_w];
assign c833ibus[temp_w*4 +:temp_w] = v1076obus[temp_w*3 +:temp_w];
assign v1076ibus[data_w*3 +:data_w] = c833obus[data_w*4 +:data_w];
assign c833ibus[temp_w*5 +:temp_w] = v1985obus[temp_w*1 +:temp_w];
assign v1985ibus[data_w*1 +:data_w] = c833obus[data_w*5 +:data_w];
assign c833ibus[temp_w*6 +:temp_w] = v2081obus[temp_w*0 +:temp_w];
assign v2081ibus[data_w*0 +:data_w] = c833obus[data_w*6 +:data_w];
assign c834ibus[temp_w*0 +:temp_w] = v78obus[temp_w*1 +:temp_w];
assign v78ibus[data_w*1 +:data_w] = c834obus[data_w*0 +:data_w];
assign c834ibus[temp_w*1 +:temp_w] = v437obus[temp_w*2 +:temp_w];
assign v437ibus[data_w*2 +:data_w] = c834obus[data_w*1 +:data_w];
assign c834ibus[temp_w*2 +:temp_w] = v570obus[temp_w*3 +:temp_w];
assign v570ibus[data_w*3 +:data_w] = c834obus[data_w*2 +:data_w];
assign c834ibus[temp_w*3 +:temp_w] = v685obus[temp_w*3 +:temp_w];
assign v685ibus[data_w*3 +:data_w] = c834obus[data_w*3 +:data_w];
assign c834ibus[temp_w*4 +:temp_w] = v1077obus[temp_w*3 +:temp_w];
assign v1077ibus[data_w*3 +:data_w] = c834obus[data_w*4 +:data_w];
assign c834ibus[temp_w*5 +:temp_w] = v1986obus[temp_w*1 +:temp_w];
assign v1986ibus[data_w*1 +:data_w] = c834obus[data_w*5 +:data_w];
assign c834ibus[temp_w*6 +:temp_w] = v2082obus[temp_w*0 +:temp_w];
assign v2082ibus[data_w*0 +:data_w] = c834obus[data_w*6 +:data_w];
assign c835ibus[temp_w*0 +:temp_w] = v79obus[temp_w*1 +:temp_w];
assign v79ibus[data_w*1 +:data_w] = c835obus[data_w*0 +:data_w];
assign c835ibus[temp_w*1 +:temp_w] = v438obus[temp_w*2 +:temp_w];
assign v438ibus[data_w*2 +:data_w] = c835obus[data_w*1 +:data_w];
assign c835ibus[temp_w*2 +:temp_w] = v571obus[temp_w*3 +:temp_w];
assign v571ibus[data_w*3 +:data_w] = c835obus[data_w*2 +:data_w];
assign c835ibus[temp_w*3 +:temp_w] = v686obus[temp_w*3 +:temp_w];
assign v686ibus[data_w*3 +:data_w] = c835obus[data_w*3 +:data_w];
assign c835ibus[temp_w*4 +:temp_w] = v1078obus[temp_w*3 +:temp_w];
assign v1078ibus[data_w*3 +:data_w] = c835obus[data_w*4 +:data_w];
assign c835ibus[temp_w*5 +:temp_w] = v1987obus[temp_w*1 +:temp_w];
assign v1987ibus[data_w*1 +:data_w] = c835obus[data_w*5 +:data_w];
assign c835ibus[temp_w*6 +:temp_w] = v2083obus[temp_w*0 +:temp_w];
assign v2083ibus[data_w*0 +:data_w] = c835obus[data_w*6 +:data_w];
assign c836ibus[temp_w*0 +:temp_w] = v80obus[temp_w*1 +:temp_w];
assign v80ibus[data_w*1 +:data_w] = c836obus[data_w*0 +:data_w];
assign c836ibus[temp_w*1 +:temp_w] = v439obus[temp_w*2 +:temp_w];
assign v439ibus[data_w*2 +:data_w] = c836obus[data_w*1 +:data_w];
assign c836ibus[temp_w*2 +:temp_w] = v572obus[temp_w*3 +:temp_w];
assign v572ibus[data_w*3 +:data_w] = c836obus[data_w*2 +:data_w];
assign c836ibus[temp_w*3 +:temp_w] = v687obus[temp_w*3 +:temp_w];
assign v687ibus[data_w*3 +:data_w] = c836obus[data_w*3 +:data_w];
assign c836ibus[temp_w*4 +:temp_w] = v1079obus[temp_w*3 +:temp_w];
assign v1079ibus[data_w*3 +:data_w] = c836obus[data_w*4 +:data_w];
assign c836ibus[temp_w*5 +:temp_w] = v1988obus[temp_w*1 +:temp_w];
assign v1988ibus[data_w*1 +:data_w] = c836obus[data_w*5 +:data_w];
assign c836ibus[temp_w*6 +:temp_w] = v2084obus[temp_w*0 +:temp_w];
assign v2084ibus[data_w*0 +:data_w] = c836obus[data_w*6 +:data_w];
assign c837ibus[temp_w*0 +:temp_w] = v81obus[temp_w*1 +:temp_w];
assign v81ibus[data_w*1 +:data_w] = c837obus[data_w*0 +:data_w];
assign c837ibus[temp_w*1 +:temp_w] = v440obus[temp_w*2 +:temp_w];
assign v440ibus[data_w*2 +:data_w] = c837obus[data_w*1 +:data_w];
assign c837ibus[temp_w*2 +:temp_w] = v573obus[temp_w*3 +:temp_w];
assign v573ibus[data_w*3 +:data_w] = c837obus[data_w*2 +:data_w];
assign c837ibus[temp_w*3 +:temp_w] = v688obus[temp_w*3 +:temp_w];
assign v688ibus[data_w*3 +:data_w] = c837obus[data_w*3 +:data_w];
assign c837ibus[temp_w*4 +:temp_w] = v1080obus[temp_w*3 +:temp_w];
assign v1080ibus[data_w*3 +:data_w] = c837obus[data_w*4 +:data_w];
assign c837ibus[temp_w*5 +:temp_w] = v1989obus[temp_w*1 +:temp_w];
assign v1989ibus[data_w*1 +:data_w] = c837obus[data_w*5 +:data_w];
assign c837ibus[temp_w*6 +:temp_w] = v2085obus[temp_w*0 +:temp_w];
assign v2085ibus[data_w*0 +:data_w] = c837obus[data_w*6 +:data_w];
assign c838ibus[temp_w*0 +:temp_w] = v82obus[temp_w*1 +:temp_w];
assign v82ibus[data_w*1 +:data_w] = c838obus[data_w*0 +:data_w];
assign c838ibus[temp_w*1 +:temp_w] = v441obus[temp_w*2 +:temp_w];
assign v441ibus[data_w*2 +:data_w] = c838obus[data_w*1 +:data_w];
assign c838ibus[temp_w*2 +:temp_w] = v574obus[temp_w*3 +:temp_w];
assign v574ibus[data_w*3 +:data_w] = c838obus[data_w*2 +:data_w];
assign c838ibus[temp_w*3 +:temp_w] = v689obus[temp_w*3 +:temp_w];
assign v689ibus[data_w*3 +:data_w] = c838obus[data_w*3 +:data_w];
assign c838ibus[temp_w*4 +:temp_w] = v1081obus[temp_w*3 +:temp_w];
assign v1081ibus[data_w*3 +:data_w] = c838obus[data_w*4 +:data_w];
assign c838ibus[temp_w*5 +:temp_w] = v1990obus[temp_w*1 +:temp_w];
assign v1990ibus[data_w*1 +:data_w] = c838obus[data_w*5 +:data_w];
assign c838ibus[temp_w*6 +:temp_w] = v2086obus[temp_w*0 +:temp_w];
assign v2086ibus[data_w*0 +:data_w] = c838obus[data_w*6 +:data_w];
assign c839ibus[temp_w*0 +:temp_w] = v83obus[temp_w*1 +:temp_w];
assign v83ibus[data_w*1 +:data_w] = c839obus[data_w*0 +:data_w];
assign c839ibus[temp_w*1 +:temp_w] = v442obus[temp_w*2 +:temp_w];
assign v442ibus[data_w*2 +:data_w] = c839obus[data_w*1 +:data_w];
assign c839ibus[temp_w*2 +:temp_w] = v575obus[temp_w*3 +:temp_w];
assign v575ibus[data_w*3 +:data_w] = c839obus[data_w*2 +:data_w];
assign c839ibus[temp_w*3 +:temp_w] = v690obus[temp_w*3 +:temp_w];
assign v690ibus[data_w*3 +:data_w] = c839obus[data_w*3 +:data_w];
assign c839ibus[temp_w*4 +:temp_w] = v1082obus[temp_w*3 +:temp_w];
assign v1082ibus[data_w*3 +:data_w] = c839obus[data_w*4 +:data_w];
assign c839ibus[temp_w*5 +:temp_w] = v1991obus[temp_w*1 +:temp_w];
assign v1991ibus[data_w*1 +:data_w] = c839obus[data_w*5 +:data_w];
assign c839ibus[temp_w*6 +:temp_w] = v2087obus[temp_w*0 +:temp_w];
assign v2087ibus[data_w*0 +:data_w] = c839obus[data_w*6 +:data_w];
assign c840ibus[temp_w*0 +:temp_w] = v84obus[temp_w*1 +:temp_w];
assign v84ibus[data_w*1 +:data_w] = c840obus[data_w*0 +:data_w];
assign c840ibus[temp_w*1 +:temp_w] = v443obus[temp_w*2 +:temp_w];
assign v443ibus[data_w*2 +:data_w] = c840obus[data_w*1 +:data_w];
assign c840ibus[temp_w*2 +:temp_w] = v480obus[temp_w*3 +:temp_w];
assign v480ibus[data_w*3 +:data_w] = c840obus[data_w*2 +:data_w];
assign c840ibus[temp_w*3 +:temp_w] = v691obus[temp_w*3 +:temp_w];
assign v691ibus[data_w*3 +:data_w] = c840obus[data_w*3 +:data_w];
assign c840ibus[temp_w*4 +:temp_w] = v1083obus[temp_w*3 +:temp_w];
assign v1083ibus[data_w*3 +:data_w] = c840obus[data_w*4 +:data_w];
assign c840ibus[temp_w*5 +:temp_w] = v1992obus[temp_w*1 +:temp_w];
assign v1992ibus[data_w*1 +:data_w] = c840obus[data_w*5 +:data_w];
assign c840ibus[temp_w*6 +:temp_w] = v2088obus[temp_w*0 +:temp_w];
assign v2088ibus[data_w*0 +:data_w] = c840obus[data_w*6 +:data_w];
assign c841ibus[temp_w*0 +:temp_w] = v85obus[temp_w*1 +:temp_w];
assign v85ibus[data_w*1 +:data_w] = c841obus[data_w*0 +:data_w];
assign c841ibus[temp_w*1 +:temp_w] = v444obus[temp_w*2 +:temp_w];
assign v444ibus[data_w*2 +:data_w] = c841obus[data_w*1 +:data_w];
assign c841ibus[temp_w*2 +:temp_w] = v481obus[temp_w*3 +:temp_w];
assign v481ibus[data_w*3 +:data_w] = c841obus[data_w*2 +:data_w];
assign c841ibus[temp_w*3 +:temp_w] = v692obus[temp_w*3 +:temp_w];
assign v692ibus[data_w*3 +:data_w] = c841obus[data_w*3 +:data_w];
assign c841ibus[temp_w*4 +:temp_w] = v1084obus[temp_w*3 +:temp_w];
assign v1084ibus[data_w*3 +:data_w] = c841obus[data_w*4 +:data_w];
assign c841ibus[temp_w*5 +:temp_w] = v1993obus[temp_w*1 +:temp_w];
assign v1993ibus[data_w*1 +:data_w] = c841obus[data_w*5 +:data_w];
assign c841ibus[temp_w*6 +:temp_w] = v2089obus[temp_w*0 +:temp_w];
assign v2089ibus[data_w*0 +:data_w] = c841obus[data_w*6 +:data_w];
assign c842ibus[temp_w*0 +:temp_w] = v86obus[temp_w*1 +:temp_w];
assign v86ibus[data_w*1 +:data_w] = c842obus[data_w*0 +:data_w];
assign c842ibus[temp_w*1 +:temp_w] = v445obus[temp_w*2 +:temp_w];
assign v445ibus[data_w*2 +:data_w] = c842obus[data_w*1 +:data_w];
assign c842ibus[temp_w*2 +:temp_w] = v482obus[temp_w*3 +:temp_w];
assign v482ibus[data_w*3 +:data_w] = c842obus[data_w*2 +:data_w];
assign c842ibus[temp_w*3 +:temp_w] = v693obus[temp_w*3 +:temp_w];
assign v693ibus[data_w*3 +:data_w] = c842obus[data_w*3 +:data_w];
assign c842ibus[temp_w*4 +:temp_w] = v1085obus[temp_w*3 +:temp_w];
assign v1085ibus[data_w*3 +:data_w] = c842obus[data_w*4 +:data_w];
assign c842ibus[temp_w*5 +:temp_w] = v1994obus[temp_w*1 +:temp_w];
assign v1994ibus[data_w*1 +:data_w] = c842obus[data_w*5 +:data_w];
assign c842ibus[temp_w*6 +:temp_w] = v2090obus[temp_w*0 +:temp_w];
assign v2090ibus[data_w*0 +:data_w] = c842obus[data_w*6 +:data_w];
assign c843ibus[temp_w*0 +:temp_w] = v87obus[temp_w*1 +:temp_w];
assign v87ibus[data_w*1 +:data_w] = c843obus[data_w*0 +:data_w];
assign c843ibus[temp_w*1 +:temp_w] = v446obus[temp_w*2 +:temp_w];
assign v446ibus[data_w*2 +:data_w] = c843obus[data_w*1 +:data_w];
assign c843ibus[temp_w*2 +:temp_w] = v483obus[temp_w*3 +:temp_w];
assign v483ibus[data_w*3 +:data_w] = c843obus[data_w*2 +:data_w];
assign c843ibus[temp_w*3 +:temp_w] = v694obus[temp_w*3 +:temp_w];
assign v694ibus[data_w*3 +:data_w] = c843obus[data_w*3 +:data_w];
assign c843ibus[temp_w*4 +:temp_w] = v1086obus[temp_w*3 +:temp_w];
assign v1086ibus[data_w*3 +:data_w] = c843obus[data_w*4 +:data_w];
assign c843ibus[temp_w*5 +:temp_w] = v1995obus[temp_w*1 +:temp_w];
assign v1995ibus[data_w*1 +:data_w] = c843obus[data_w*5 +:data_w];
assign c843ibus[temp_w*6 +:temp_w] = v2091obus[temp_w*0 +:temp_w];
assign v2091ibus[data_w*0 +:data_w] = c843obus[data_w*6 +:data_w];
assign c844ibus[temp_w*0 +:temp_w] = v88obus[temp_w*1 +:temp_w];
assign v88ibus[data_w*1 +:data_w] = c844obus[data_w*0 +:data_w];
assign c844ibus[temp_w*1 +:temp_w] = v447obus[temp_w*2 +:temp_w];
assign v447ibus[data_w*2 +:data_w] = c844obus[data_w*1 +:data_w];
assign c844ibus[temp_w*2 +:temp_w] = v484obus[temp_w*3 +:temp_w];
assign v484ibus[data_w*3 +:data_w] = c844obus[data_w*2 +:data_w];
assign c844ibus[temp_w*3 +:temp_w] = v695obus[temp_w*3 +:temp_w];
assign v695ibus[data_w*3 +:data_w] = c844obus[data_w*3 +:data_w];
assign c844ibus[temp_w*4 +:temp_w] = v1087obus[temp_w*3 +:temp_w];
assign v1087ibus[data_w*3 +:data_w] = c844obus[data_w*4 +:data_w];
assign c844ibus[temp_w*5 +:temp_w] = v1996obus[temp_w*1 +:temp_w];
assign v1996ibus[data_w*1 +:data_w] = c844obus[data_w*5 +:data_w];
assign c844ibus[temp_w*6 +:temp_w] = v2092obus[temp_w*0 +:temp_w];
assign v2092ibus[data_w*0 +:data_w] = c844obus[data_w*6 +:data_w];
assign c845ibus[temp_w*0 +:temp_w] = v89obus[temp_w*1 +:temp_w];
assign v89ibus[data_w*1 +:data_w] = c845obus[data_w*0 +:data_w];
assign c845ibus[temp_w*1 +:temp_w] = v448obus[temp_w*2 +:temp_w];
assign v448ibus[data_w*2 +:data_w] = c845obus[data_w*1 +:data_w];
assign c845ibus[temp_w*2 +:temp_w] = v485obus[temp_w*3 +:temp_w];
assign v485ibus[data_w*3 +:data_w] = c845obus[data_w*2 +:data_w];
assign c845ibus[temp_w*3 +:temp_w] = v696obus[temp_w*3 +:temp_w];
assign v696ibus[data_w*3 +:data_w] = c845obus[data_w*3 +:data_w];
assign c845ibus[temp_w*4 +:temp_w] = v1088obus[temp_w*3 +:temp_w];
assign v1088ibus[data_w*3 +:data_w] = c845obus[data_w*4 +:data_w];
assign c845ibus[temp_w*5 +:temp_w] = v1997obus[temp_w*1 +:temp_w];
assign v1997ibus[data_w*1 +:data_w] = c845obus[data_w*5 +:data_w];
assign c845ibus[temp_w*6 +:temp_w] = v2093obus[temp_w*0 +:temp_w];
assign v2093ibus[data_w*0 +:data_w] = c845obus[data_w*6 +:data_w];
assign c846ibus[temp_w*0 +:temp_w] = v90obus[temp_w*1 +:temp_w];
assign v90ibus[data_w*1 +:data_w] = c846obus[data_w*0 +:data_w];
assign c846ibus[temp_w*1 +:temp_w] = v449obus[temp_w*2 +:temp_w];
assign v449ibus[data_w*2 +:data_w] = c846obus[data_w*1 +:data_w];
assign c846ibus[temp_w*2 +:temp_w] = v486obus[temp_w*3 +:temp_w];
assign v486ibus[data_w*3 +:data_w] = c846obus[data_w*2 +:data_w];
assign c846ibus[temp_w*3 +:temp_w] = v697obus[temp_w*3 +:temp_w];
assign v697ibus[data_w*3 +:data_w] = c846obus[data_w*3 +:data_w];
assign c846ibus[temp_w*4 +:temp_w] = v1089obus[temp_w*3 +:temp_w];
assign v1089ibus[data_w*3 +:data_w] = c846obus[data_w*4 +:data_w];
assign c846ibus[temp_w*5 +:temp_w] = v1998obus[temp_w*1 +:temp_w];
assign v1998ibus[data_w*1 +:data_w] = c846obus[data_w*5 +:data_w];
assign c846ibus[temp_w*6 +:temp_w] = v2094obus[temp_w*0 +:temp_w];
assign v2094ibus[data_w*0 +:data_w] = c846obus[data_w*6 +:data_w];
assign c847ibus[temp_w*0 +:temp_w] = v91obus[temp_w*1 +:temp_w];
assign v91ibus[data_w*1 +:data_w] = c847obus[data_w*0 +:data_w];
assign c847ibus[temp_w*1 +:temp_w] = v450obus[temp_w*2 +:temp_w];
assign v450ibus[data_w*2 +:data_w] = c847obus[data_w*1 +:data_w];
assign c847ibus[temp_w*2 +:temp_w] = v487obus[temp_w*3 +:temp_w];
assign v487ibus[data_w*3 +:data_w] = c847obus[data_w*2 +:data_w];
assign c847ibus[temp_w*3 +:temp_w] = v698obus[temp_w*3 +:temp_w];
assign v698ibus[data_w*3 +:data_w] = c847obus[data_w*3 +:data_w];
assign c847ibus[temp_w*4 +:temp_w] = v1090obus[temp_w*3 +:temp_w];
assign v1090ibus[data_w*3 +:data_w] = c847obus[data_w*4 +:data_w];
assign c847ibus[temp_w*5 +:temp_w] = v1999obus[temp_w*1 +:temp_w];
assign v1999ibus[data_w*1 +:data_w] = c847obus[data_w*5 +:data_w];
assign c847ibus[temp_w*6 +:temp_w] = v2095obus[temp_w*0 +:temp_w];
assign v2095ibus[data_w*0 +:data_w] = c847obus[data_w*6 +:data_w];
assign c848ibus[temp_w*0 +:temp_w] = v92obus[temp_w*1 +:temp_w];
assign v92ibus[data_w*1 +:data_w] = c848obus[data_w*0 +:data_w];
assign c848ibus[temp_w*1 +:temp_w] = v451obus[temp_w*2 +:temp_w];
assign v451ibus[data_w*2 +:data_w] = c848obus[data_w*1 +:data_w];
assign c848ibus[temp_w*2 +:temp_w] = v488obus[temp_w*3 +:temp_w];
assign v488ibus[data_w*3 +:data_w] = c848obus[data_w*2 +:data_w];
assign c848ibus[temp_w*3 +:temp_w] = v699obus[temp_w*3 +:temp_w];
assign v699ibus[data_w*3 +:data_w] = c848obus[data_w*3 +:data_w];
assign c848ibus[temp_w*4 +:temp_w] = v1091obus[temp_w*3 +:temp_w];
assign v1091ibus[data_w*3 +:data_w] = c848obus[data_w*4 +:data_w];
assign c848ibus[temp_w*5 +:temp_w] = v2000obus[temp_w*1 +:temp_w];
assign v2000ibus[data_w*1 +:data_w] = c848obus[data_w*5 +:data_w];
assign c848ibus[temp_w*6 +:temp_w] = v2096obus[temp_w*0 +:temp_w];
assign v2096ibus[data_w*0 +:data_w] = c848obus[data_w*6 +:data_w];
assign c849ibus[temp_w*0 +:temp_w] = v93obus[temp_w*1 +:temp_w];
assign v93ibus[data_w*1 +:data_w] = c849obus[data_w*0 +:data_w];
assign c849ibus[temp_w*1 +:temp_w] = v452obus[temp_w*2 +:temp_w];
assign v452ibus[data_w*2 +:data_w] = c849obus[data_w*1 +:data_w];
assign c849ibus[temp_w*2 +:temp_w] = v489obus[temp_w*3 +:temp_w];
assign v489ibus[data_w*3 +:data_w] = c849obus[data_w*2 +:data_w];
assign c849ibus[temp_w*3 +:temp_w] = v700obus[temp_w*3 +:temp_w];
assign v700ibus[data_w*3 +:data_w] = c849obus[data_w*3 +:data_w];
assign c849ibus[temp_w*4 +:temp_w] = v1092obus[temp_w*3 +:temp_w];
assign v1092ibus[data_w*3 +:data_w] = c849obus[data_w*4 +:data_w];
assign c849ibus[temp_w*5 +:temp_w] = v2001obus[temp_w*1 +:temp_w];
assign v2001ibus[data_w*1 +:data_w] = c849obus[data_w*5 +:data_w];
assign c849ibus[temp_w*6 +:temp_w] = v2097obus[temp_w*0 +:temp_w];
assign v2097ibus[data_w*0 +:data_w] = c849obus[data_w*6 +:data_w];
assign c850ibus[temp_w*0 +:temp_w] = v94obus[temp_w*1 +:temp_w];
assign v94ibus[data_w*1 +:data_w] = c850obus[data_w*0 +:data_w];
assign c850ibus[temp_w*1 +:temp_w] = v453obus[temp_w*2 +:temp_w];
assign v453ibus[data_w*2 +:data_w] = c850obus[data_w*1 +:data_w];
assign c850ibus[temp_w*2 +:temp_w] = v490obus[temp_w*3 +:temp_w];
assign v490ibus[data_w*3 +:data_w] = c850obus[data_w*2 +:data_w];
assign c850ibus[temp_w*3 +:temp_w] = v701obus[temp_w*3 +:temp_w];
assign v701ibus[data_w*3 +:data_w] = c850obus[data_w*3 +:data_w];
assign c850ibus[temp_w*4 +:temp_w] = v1093obus[temp_w*3 +:temp_w];
assign v1093ibus[data_w*3 +:data_w] = c850obus[data_w*4 +:data_w];
assign c850ibus[temp_w*5 +:temp_w] = v2002obus[temp_w*1 +:temp_w];
assign v2002ibus[data_w*1 +:data_w] = c850obus[data_w*5 +:data_w];
assign c850ibus[temp_w*6 +:temp_w] = v2098obus[temp_w*0 +:temp_w];
assign v2098ibus[data_w*0 +:data_w] = c850obus[data_w*6 +:data_w];
assign c851ibus[temp_w*0 +:temp_w] = v95obus[temp_w*1 +:temp_w];
assign v95ibus[data_w*1 +:data_w] = c851obus[data_w*0 +:data_w];
assign c851ibus[temp_w*1 +:temp_w] = v454obus[temp_w*2 +:temp_w];
assign v454ibus[data_w*2 +:data_w] = c851obus[data_w*1 +:data_w];
assign c851ibus[temp_w*2 +:temp_w] = v491obus[temp_w*3 +:temp_w];
assign v491ibus[data_w*3 +:data_w] = c851obus[data_w*2 +:data_w];
assign c851ibus[temp_w*3 +:temp_w] = v702obus[temp_w*3 +:temp_w];
assign v702ibus[data_w*3 +:data_w] = c851obus[data_w*3 +:data_w];
assign c851ibus[temp_w*4 +:temp_w] = v1094obus[temp_w*3 +:temp_w];
assign v1094ibus[data_w*3 +:data_w] = c851obus[data_w*4 +:data_w];
assign c851ibus[temp_w*5 +:temp_w] = v2003obus[temp_w*1 +:temp_w];
assign v2003ibus[data_w*1 +:data_w] = c851obus[data_w*5 +:data_w];
assign c851ibus[temp_w*6 +:temp_w] = v2099obus[temp_w*0 +:temp_w];
assign v2099ibus[data_w*0 +:data_w] = c851obus[data_w*6 +:data_w];
assign c852ibus[temp_w*0 +:temp_w] = v0obus[temp_w*1 +:temp_w];
assign v0ibus[data_w*1 +:data_w] = c852obus[data_w*0 +:data_w];
assign c852ibus[temp_w*1 +:temp_w] = v455obus[temp_w*2 +:temp_w];
assign v455ibus[data_w*2 +:data_w] = c852obus[data_w*1 +:data_w];
assign c852ibus[temp_w*2 +:temp_w] = v492obus[temp_w*3 +:temp_w];
assign v492ibus[data_w*3 +:data_w] = c852obus[data_w*2 +:data_w];
assign c852ibus[temp_w*3 +:temp_w] = v703obus[temp_w*3 +:temp_w];
assign v703ibus[data_w*3 +:data_w] = c852obus[data_w*3 +:data_w];
assign c852ibus[temp_w*4 +:temp_w] = v1095obus[temp_w*3 +:temp_w];
assign v1095ibus[data_w*3 +:data_w] = c852obus[data_w*4 +:data_w];
assign c852ibus[temp_w*5 +:temp_w] = v2004obus[temp_w*1 +:temp_w];
assign v2004ibus[data_w*1 +:data_w] = c852obus[data_w*5 +:data_w];
assign c852ibus[temp_w*6 +:temp_w] = v2100obus[temp_w*0 +:temp_w];
assign v2100ibus[data_w*0 +:data_w] = c852obus[data_w*6 +:data_w];
assign c853ibus[temp_w*0 +:temp_w] = v1obus[temp_w*1 +:temp_w];
assign v1ibus[data_w*1 +:data_w] = c853obus[data_w*0 +:data_w];
assign c853ibus[temp_w*1 +:temp_w] = v456obus[temp_w*2 +:temp_w];
assign v456ibus[data_w*2 +:data_w] = c853obus[data_w*1 +:data_w];
assign c853ibus[temp_w*2 +:temp_w] = v493obus[temp_w*3 +:temp_w];
assign v493ibus[data_w*3 +:data_w] = c853obus[data_w*2 +:data_w];
assign c853ibus[temp_w*3 +:temp_w] = v704obus[temp_w*3 +:temp_w];
assign v704ibus[data_w*3 +:data_w] = c853obus[data_w*3 +:data_w];
assign c853ibus[temp_w*4 +:temp_w] = v1096obus[temp_w*3 +:temp_w];
assign v1096ibus[data_w*3 +:data_w] = c853obus[data_w*4 +:data_w];
assign c853ibus[temp_w*5 +:temp_w] = v2005obus[temp_w*1 +:temp_w];
assign v2005ibus[data_w*1 +:data_w] = c853obus[data_w*5 +:data_w];
assign c853ibus[temp_w*6 +:temp_w] = v2101obus[temp_w*0 +:temp_w];
assign v2101ibus[data_w*0 +:data_w] = c853obus[data_w*6 +:data_w];
assign c854ibus[temp_w*0 +:temp_w] = v2obus[temp_w*1 +:temp_w];
assign v2ibus[data_w*1 +:data_w] = c854obus[data_w*0 +:data_w];
assign c854ibus[temp_w*1 +:temp_w] = v457obus[temp_w*2 +:temp_w];
assign v457ibus[data_w*2 +:data_w] = c854obus[data_w*1 +:data_w];
assign c854ibus[temp_w*2 +:temp_w] = v494obus[temp_w*3 +:temp_w];
assign v494ibus[data_w*3 +:data_w] = c854obus[data_w*2 +:data_w];
assign c854ibus[temp_w*3 +:temp_w] = v705obus[temp_w*3 +:temp_w];
assign v705ibus[data_w*3 +:data_w] = c854obus[data_w*3 +:data_w];
assign c854ibus[temp_w*4 +:temp_w] = v1097obus[temp_w*3 +:temp_w];
assign v1097ibus[data_w*3 +:data_w] = c854obus[data_w*4 +:data_w];
assign c854ibus[temp_w*5 +:temp_w] = v2006obus[temp_w*1 +:temp_w];
assign v2006ibus[data_w*1 +:data_w] = c854obus[data_w*5 +:data_w];
assign c854ibus[temp_w*6 +:temp_w] = v2102obus[temp_w*0 +:temp_w];
assign v2102ibus[data_w*0 +:data_w] = c854obus[data_w*6 +:data_w];
assign c855ibus[temp_w*0 +:temp_w] = v3obus[temp_w*1 +:temp_w];
assign v3ibus[data_w*1 +:data_w] = c855obus[data_w*0 +:data_w];
assign c855ibus[temp_w*1 +:temp_w] = v458obus[temp_w*2 +:temp_w];
assign v458ibus[data_w*2 +:data_w] = c855obus[data_w*1 +:data_w];
assign c855ibus[temp_w*2 +:temp_w] = v495obus[temp_w*3 +:temp_w];
assign v495ibus[data_w*3 +:data_w] = c855obus[data_w*2 +:data_w];
assign c855ibus[temp_w*3 +:temp_w] = v706obus[temp_w*3 +:temp_w];
assign v706ibus[data_w*3 +:data_w] = c855obus[data_w*3 +:data_w];
assign c855ibus[temp_w*4 +:temp_w] = v1098obus[temp_w*3 +:temp_w];
assign v1098ibus[data_w*3 +:data_w] = c855obus[data_w*4 +:data_w];
assign c855ibus[temp_w*5 +:temp_w] = v2007obus[temp_w*1 +:temp_w];
assign v2007ibus[data_w*1 +:data_w] = c855obus[data_w*5 +:data_w];
assign c855ibus[temp_w*6 +:temp_w] = v2103obus[temp_w*0 +:temp_w];
assign v2103ibus[data_w*0 +:data_w] = c855obus[data_w*6 +:data_w];
assign c856ibus[temp_w*0 +:temp_w] = v4obus[temp_w*1 +:temp_w];
assign v4ibus[data_w*1 +:data_w] = c856obus[data_w*0 +:data_w];
assign c856ibus[temp_w*1 +:temp_w] = v459obus[temp_w*2 +:temp_w];
assign v459ibus[data_w*2 +:data_w] = c856obus[data_w*1 +:data_w];
assign c856ibus[temp_w*2 +:temp_w] = v496obus[temp_w*3 +:temp_w];
assign v496ibus[data_w*3 +:data_w] = c856obus[data_w*2 +:data_w];
assign c856ibus[temp_w*3 +:temp_w] = v707obus[temp_w*3 +:temp_w];
assign v707ibus[data_w*3 +:data_w] = c856obus[data_w*3 +:data_w];
assign c856ibus[temp_w*4 +:temp_w] = v1099obus[temp_w*3 +:temp_w];
assign v1099ibus[data_w*3 +:data_w] = c856obus[data_w*4 +:data_w];
assign c856ibus[temp_w*5 +:temp_w] = v2008obus[temp_w*1 +:temp_w];
assign v2008ibus[data_w*1 +:data_w] = c856obus[data_w*5 +:data_w];
assign c856ibus[temp_w*6 +:temp_w] = v2104obus[temp_w*0 +:temp_w];
assign v2104ibus[data_w*0 +:data_w] = c856obus[data_w*6 +:data_w];
assign c857ibus[temp_w*0 +:temp_w] = v5obus[temp_w*1 +:temp_w];
assign v5ibus[data_w*1 +:data_w] = c857obus[data_w*0 +:data_w];
assign c857ibus[temp_w*1 +:temp_w] = v460obus[temp_w*2 +:temp_w];
assign v460ibus[data_w*2 +:data_w] = c857obus[data_w*1 +:data_w];
assign c857ibus[temp_w*2 +:temp_w] = v497obus[temp_w*3 +:temp_w];
assign v497ibus[data_w*3 +:data_w] = c857obus[data_w*2 +:data_w];
assign c857ibus[temp_w*3 +:temp_w] = v708obus[temp_w*3 +:temp_w];
assign v708ibus[data_w*3 +:data_w] = c857obus[data_w*3 +:data_w];
assign c857ibus[temp_w*4 +:temp_w] = v1100obus[temp_w*3 +:temp_w];
assign v1100ibus[data_w*3 +:data_w] = c857obus[data_w*4 +:data_w];
assign c857ibus[temp_w*5 +:temp_w] = v2009obus[temp_w*1 +:temp_w];
assign v2009ibus[data_w*1 +:data_w] = c857obus[data_w*5 +:data_w];
assign c857ibus[temp_w*6 +:temp_w] = v2105obus[temp_w*0 +:temp_w];
assign v2105ibus[data_w*0 +:data_w] = c857obus[data_w*6 +:data_w];
assign c858ibus[temp_w*0 +:temp_w] = v6obus[temp_w*1 +:temp_w];
assign v6ibus[data_w*1 +:data_w] = c858obus[data_w*0 +:data_w];
assign c858ibus[temp_w*1 +:temp_w] = v461obus[temp_w*2 +:temp_w];
assign v461ibus[data_w*2 +:data_w] = c858obus[data_w*1 +:data_w];
assign c858ibus[temp_w*2 +:temp_w] = v498obus[temp_w*3 +:temp_w];
assign v498ibus[data_w*3 +:data_w] = c858obus[data_w*2 +:data_w];
assign c858ibus[temp_w*3 +:temp_w] = v709obus[temp_w*3 +:temp_w];
assign v709ibus[data_w*3 +:data_w] = c858obus[data_w*3 +:data_w];
assign c858ibus[temp_w*4 +:temp_w] = v1101obus[temp_w*3 +:temp_w];
assign v1101ibus[data_w*3 +:data_w] = c858obus[data_w*4 +:data_w];
assign c858ibus[temp_w*5 +:temp_w] = v2010obus[temp_w*1 +:temp_w];
assign v2010ibus[data_w*1 +:data_w] = c858obus[data_w*5 +:data_w];
assign c858ibus[temp_w*6 +:temp_w] = v2106obus[temp_w*0 +:temp_w];
assign v2106ibus[data_w*0 +:data_w] = c858obus[data_w*6 +:data_w];
assign c859ibus[temp_w*0 +:temp_w] = v7obus[temp_w*1 +:temp_w];
assign v7ibus[data_w*1 +:data_w] = c859obus[data_w*0 +:data_w];
assign c859ibus[temp_w*1 +:temp_w] = v462obus[temp_w*2 +:temp_w];
assign v462ibus[data_w*2 +:data_w] = c859obus[data_w*1 +:data_w];
assign c859ibus[temp_w*2 +:temp_w] = v499obus[temp_w*3 +:temp_w];
assign v499ibus[data_w*3 +:data_w] = c859obus[data_w*2 +:data_w];
assign c859ibus[temp_w*3 +:temp_w] = v710obus[temp_w*3 +:temp_w];
assign v710ibus[data_w*3 +:data_w] = c859obus[data_w*3 +:data_w];
assign c859ibus[temp_w*4 +:temp_w] = v1102obus[temp_w*3 +:temp_w];
assign v1102ibus[data_w*3 +:data_w] = c859obus[data_w*4 +:data_w];
assign c859ibus[temp_w*5 +:temp_w] = v2011obus[temp_w*1 +:temp_w];
assign v2011ibus[data_w*1 +:data_w] = c859obus[data_w*5 +:data_w];
assign c859ibus[temp_w*6 +:temp_w] = v2107obus[temp_w*0 +:temp_w];
assign v2107ibus[data_w*0 +:data_w] = c859obus[data_w*6 +:data_w];
assign c860ibus[temp_w*0 +:temp_w] = v8obus[temp_w*1 +:temp_w];
assign v8ibus[data_w*1 +:data_w] = c860obus[data_w*0 +:data_w];
assign c860ibus[temp_w*1 +:temp_w] = v463obus[temp_w*2 +:temp_w];
assign v463ibus[data_w*2 +:data_w] = c860obus[data_w*1 +:data_w];
assign c860ibus[temp_w*2 +:temp_w] = v500obus[temp_w*3 +:temp_w];
assign v500ibus[data_w*3 +:data_w] = c860obus[data_w*2 +:data_w];
assign c860ibus[temp_w*3 +:temp_w] = v711obus[temp_w*3 +:temp_w];
assign v711ibus[data_w*3 +:data_w] = c860obus[data_w*3 +:data_w];
assign c860ibus[temp_w*4 +:temp_w] = v1103obus[temp_w*3 +:temp_w];
assign v1103ibus[data_w*3 +:data_w] = c860obus[data_w*4 +:data_w];
assign c860ibus[temp_w*5 +:temp_w] = v2012obus[temp_w*1 +:temp_w];
assign v2012ibus[data_w*1 +:data_w] = c860obus[data_w*5 +:data_w];
assign c860ibus[temp_w*6 +:temp_w] = v2108obus[temp_w*0 +:temp_w];
assign v2108ibus[data_w*0 +:data_w] = c860obus[data_w*6 +:data_w];
assign c861ibus[temp_w*0 +:temp_w] = v9obus[temp_w*1 +:temp_w];
assign v9ibus[data_w*1 +:data_w] = c861obus[data_w*0 +:data_w];
assign c861ibus[temp_w*1 +:temp_w] = v464obus[temp_w*2 +:temp_w];
assign v464ibus[data_w*2 +:data_w] = c861obus[data_w*1 +:data_w];
assign c861ibus[temp_w*2 +:temp_w] = v501obus[temp_w*3 +:temp_w];
assign v501ibus[data_w*3 +:data_w] = c861obus[data_w*2 +:data_w];
assign c861ibus[temp_w*3 +:temp_w] = v712obus[temp_w*3 +:temp_w];
assign v712ibus[data_w*3 +:data_w] = c861obus[data_w*3 +:data_w];
assign c861ibus[temp_w*4 +:temp_w] = v1104obus[temp_w*3 +:temp_w];
assign v1104ibus[data_w*3 +:data_w] = c861obus[data_w*4 +:data_w];
assign c861ibus[temp_w*5 +:temp_w] = v2013obus[temp_w*1 +:temp_w];
assign v2013ibus[data_w*1 +:data_w] = c861obus[data_w*5 +:data_w];
assign c861ibus[temp_w*6 +:temp_w] = v2109obus[temp_w*0 +:temp_w];
assign v2109ibus[data_w*0 +:data_w] = c861obus[data_w*6 +:data_w];
assign c862ibus[temp_w*0 +:temp_w] = v10obus[temp_w*1 +:temp_w];
assign v10ibus[data_w*1 +:data_w] = c862obus[data_w*0 +:data_w];
assign c862ibus[temp_w*1 +:temp_w] = v465obus[temp_w*2 +:temp_w];
assign v465ibus[data_w*2 +:data_w] = c862obus[data_w*1 +:data_w];
assign c862ibus[temp_w*2 +:temp_w] = v502obus[temp_w*3 +:temp_w];
assign v502ibus[data_w*3 +:data_w] = c862obus[data_w*2 +:data_w];
assign c862ibus[temp_w*3 +:temp_w] = v713obus[temp_w*3 +:temp_w];
assign v713ibus[data_w*3 +:data_w] = c862obus[data_w*3 +:data_w];
assign c862ibus[temp_w*4 +:temp_w] = v1105obus[temp_w*3 +:temp_w];
assign v1105ibus[data_w*3 +:data_w] = c862obus[data_w*4 +:data_w];
assign c862ibus[temp_w*5 +:temp_w] = v2014obus[temp_w*1 +:temp_w];
assign v2014ibus[data_w*1 +:data_w] = c862obus[data_w*5 +:data_w];
assign c862ibus[temp_w*6 +:temp_w] = v2110obus[temp_w*0 +:temp_w];
assign v2110ibus[data_w*0 +:data_w] = c862obus[data_w*6 +:data_w];
assign c863ibus[temp_w*0 +:temp_w] = v11obus[temp_w*1 +:temp_w];
assign v11ibus[data_w*1 +:data_w] = c863obus[data_w*0 +:data_w];
assign c863ibus[temp_w*1 +:temp_w] = v466obus[temp_w*2 +:temp_w];
assign v466ibus[data_w*2 +:data_w] = c863obus[data_w*1 +:data_w];
assign c863ibus[temp_w*2 +:temp_w] = v503obus[temp_w*3 +:temp_w];
assign v503ibus[data_w*3 +:data_w] = c863obus[data_w*2 +:data_w];
assign c863ibus[temp_w*3 +:temp_w] = v714obus[temp_w*3 +:temp_w];
assign v714ibus[data_w*3 +:data_w] = c863obus[data_w*3 +:data_w];
assign c863ibus[temp_w*4 +:temp_w] = v1106obus[temp_w*3 +:temp_w];
assign v1106ibus[data_w*3 +:data_w] = c863obus[data_w*4 +:data_w];
assign c863ibus[temp_w*5 +:temp_w] = v2015obus[temp_w*1 +:temp_w];
assign v2015ibus[data_w*1 +:data_w] = c863obus[data_w*5 +:data_w];
assign c863ibus[temp_w*6 +:temp_w] = v2111obus[temp_w*0 +:temp_w];
assign v2111ibus[data_w*0 +:data_w] = c863obus[data_w*6 +:data_w];
assign c864ibus[temp_w*0 +:temp_w] = v574obus[temp_w*4 +:temp_w];
assign v574ibus[data_w*4 +:data_w] = c864obus[data_w*0 +:data_w];
assign c864ibus[temp_w*1 +:temp_w] = v731obus[temp_w*4 +:temp_w];
assign v731ibus[data_w*4 +:data_w] = c864obus[data_w*1 +:data_w];
assign c864ibus[temp_w*2 +:temp_w] = v1030obus[temp_w*2 +:temp_w];
assign v1030ibus[data_w*2 +:data_w] = c864obus[data_w*2 +:data_w];
assign c864ibus[temp_w*3 +:temp_w] = v1128obus[temp_w*4 +:temp_w];
assign v1128ibus[data_w*4 +:data_w] = c864obus[data_w*3 +:data_w];
assign c864ibus[temp_w*4 +:temp_w] = v2016obus[temp_w*1 +:temp_w];
assign v2016ibus[data_w*1 +:data_w] = c864obus[data_w*4 +:data_w];
assign c864ibus[temp_w*5 +:temp_w] = v2112obus[temp_w*0 +:temp_w];
assign v2112ibus[data_w*0 +:data_w] = c864obus[data_w*5 +:data_w];
assign c865ibus[temp_w*0 +:temp_w] = v575obus[temp_w*4 +:temp_w];
assign v575ibus[data_w*4 +:data_w] = c865obus[data_w*0 +:data_w];
assign c865ibus[temp_w*1 +:temp_w] = v732obus[temp_w*4 +:temp_w];
assign v732ibus[data_w*4 +:data_w] = c865obus[data_w*1 +:data_w];
assign c865ibus[temp_w*2 +:temp_w] = v1031obus[temp_w*2 +:temp_w];
assign v1031ibus[data_w*2 +:data_w] = c865obus[data_w*2 +:data_w];
assign c865ibus[temp_w*3 +:temp_w] = v1129obus[temp_w*4 +:temp_w];
assign v1129ibus[data_w*4 +:data_w] = c865obus[data_w*3 +:data_w];
assign c865ibus[temp_w*4 +:temp_w] = v2017obus[temp_w*1 +:temp_w];
assign v2017ibus[data_w*1 +:data_w] = c865obus[data_w*4 +:data_w];
assign c865ibus[temp_w*5 +:temp_w] = v2113obus[temp_w*0 +:temp_w];
assign v2113ibus[data_w*0 +:data_w] = c865obus[data_w*5 +:data_w];
assign c866ibus[temp_w*0 +:temp_w] = v480obus[temp_w*4 +:temp_w];
assign v480ibus[data_w*4 +:data_w] = c866obus[data_w*0 +:data_w];
assign c866ibus[temp_w*1 +:temp_w] = v733obus[temp_w*4 +:temp_w];
assign v733ibus[data_w*4 +:data_w] = c866obus[data_w*1 +:data_w];
assign c866ibus[temp_w*2 +:temp_w] = v1032obus[temp_w*2 +:temp_w];
assign v1032ibus[data_w*2 +:data_w] = c866obus[data_w*2 +:data_w];
assign c866ibus[temp_w*3 +:temp_w] = v1130obus[temp_w*4 +:temp_w];
assign v1130ibus[data_w*4 +:data_w] = c866obus[data_w*3 +:data_w];
assign c866ibus[temp_w*4 +:temp_w] = v2018obus[temp_w*1 +:temp_w];
assign v2018ibus[data_w*1 +:data_w] = c866obus[data_w*4 +:data_w];
assign c866ibus[temp_w*5 +:temp_w] = v2114obus[temp_w*0 +:temp_w];
assign v2114ibus[data_w*0 +:data_w] = c866obus[data_w*5 +:data_w];
assign c867ibus[temp_w*0 +:temp_w] = v481obus[temp_w*4 +:temp_w];
assign v481ibus[data_w*4 +:data_w] = c867obus[data_w*0 +:data_w];
assign c867ibus[temp_w*1 +:temp_w] = v734obus[temp_w*4 +:temp_w];
assign v734ibus[data_w*4 +:data_w] = c867obus[data_w*1 +:data_w];
assign c867ibus[temp_w*2 +:temp_w] = v1033obus[temp_w*2 +:temp_w];
assign v1033ibus[data_w*2 +:data_w] = c867obus[data_w*2 +:data_w];
assign c867ibus[temp_w*3 +:temp_w] = v1131obus[temp_w*4 +:temp_w];
assign v1131ibus[data_w*4 +:data_w] = c867obus[data_w*3 +:data_w];
assign c867ibus[temp_w*4 +:temp_w] = v2019obus[temp_w*1 +:temp_w];
assign v2019ibus[data_w*1 +:data_w] = c867obus[data_w*4 +:data_w];
assign c867ibus[temp_w*5 +:temp_w] = v2115obus[temp_w*0 +:temp_w];
assign v2115ibus[data_w*0 +:data_w] = c867obus[data_w*5 +:data_w];
assign c868ibus[temp_w*0 +:temp_w] = v482obus[temp_w*4 +:temp_w];
assign v482ibus[data_w*4 +:data_w] = c868obus[data_w*0 +:data_w];
assign c868ibus[temp_w*1 +:temp_w] = v735obus[temp_w*4 +:temp_w];
assign v735ibus[data_w*4 +:data_w] = c868obus[data_w*1 +:data_w];
assign c868ibus[temp_w*2 +:temp_w] = v1034obus[temp_w*2 +:temp_w];
assign v1034ibus[data_w*2 +:data_w] = c868obus[data_w*2 +:data_w];
assign c868ibus[temp_w*3 +:temp_w] = v1132obus[temp_w*4 +:temp_w];
assign v1132ibus[data_w*4 +:data_w] = c868obus[data_w*3 +:data_w];
assign c868ibus[temp_w*4 +:temp_w] = v2020obus[temp_w*1 +:temp_w];
assign v2020ibus[data_w*1 +:data_w] = c868obus[data_w*4 +:data_w];
assign c868ibus[temp_w*5 +:temp_w] = v2116obus[temp_w*0 +:temp_w];
assign v2116ibus[data_w*0 +:data_w] = c868obus[data_w*5 +:data_w];
assign c869ibus[temp_w*0 +:temp_w] = v483obus[temp_w*4 +:temp_w];
assign v483ibus[data_w*4 +:data_w] = c869obus[data_w*0 +:data_w];
assign c869ibus[temp_w*1 +:temp_w] = v736obus[temp_w*4 +:temp_w];
assign v736ibus[data_w*4 +:data_w] = c869obus[data_w*1 +:data_w];
assign c869ibus[temp_w*2 +:temp_w] = v1035obus[temp_w*2 +:temp_w];
assign v1035ibus[data_w*2 +:data_w] = c869obus[data_w*2 +:data_w];
assign c869ibus[temp_w*3 +:temp_w] = v1133obus[temp_w*4 +:temp_w];
assign v1133ibus[data_w*4 +:data_w] = c869obus[data_w*3 +:data_w];
assign c869ibus[temp_w*4 +:temp_w] = v2021obus[temp_w*1 +:temp_w];
assign v2021ibus[data_w*1 +:data_w] = c869obus[data_w*4 +:data_w];
assign c869ibus[temp_w*5 +:temp_w] = v2117obus[temp_w*0 +:temp_w];
assign v2117ibus[data_w*0 +:data_w] = c869obus[data_w*5 +:data_w];
assign c870ibus[temp_w*0 +:temp_w] = v484obus[temp_w*4 +:temp_w];
assign v484ibus[data_w*4 +:data_w] = c870obus[data_w*0 +:data_w];
assign c870ibus[temp_w*1 +:temp_w] = v737obus[temp_w*4 +:temp_w];
assign v737ibus[data_w*4 +:data_w] = c870obus[data_w*1 +:data_w];
assign c870ibus[temp_w*2 +:temp_w] = v1036obus[temp_w*2 +:temp_w];
assign v1036ibus[data_w*2 +:data_w] = c870obus[data_w*2 +:data_w];
assign c870ibus[temp_w*3 +:temp_w] = v1134obus[temp_w*4 +:temp_w];
assign v1134ibus[data_w*4 +:data_w] = c870obus[data_w*3 +:data_w];
assign c870ibus[temp_w*4 +:temp_w] = v2022obus[temp_w*1 +:temp_w];
assign v2022ibus[data_w*1 +:data_w] = c870obus[data_w*4 +:data_w];
assign c870ibus[temp_w*5 +:temp_w] = v2118obus[temp_w*0 +:temp_w];
assign v2118ibus[data_w*0 +:data_w] = c870obus[data_w*5 +:data_w];
assign c871ibus[temp_w*0 +:temp_w] = v485obus[temp_w*4 +:temp_w];
assign v485ibus[data_w*4 +:data_w] = c871obus[data_w*0 +:data_w];
assign c871ibus[temp_w*1 +:temp_w] = v738obus[temp_w*4 +:temp_w];
assign v738ibus[data_w*4 +:data_w] = c871obus[data_w*1 +:data_w];
assign c871ibus[temp_w*2 +:temp_w] = v1037obus[temp_w*2 +:temp_w];
assign v1037ibus[data_w*2 +:data_w] = c871obus[data_w*2 +:data_w];
assign c871ibus[temp_w*3 +:temp_w] = v1135obus[temp_w*4 +:temp_w];
assign v1135ibus[data_w*4 +:data_w] = c871obus[data_w*3 +:data_w];
assign c871ibus[temp_w*4 +:temp_w] = v2023obus[temp_w*1 +:temp_w];
assign v2023ibus[data_w*1 +:data_w] = c871obus[data_w*4 +:data_w];
assign c871ibus[temp_w*5 +:temp_w] = v2119obus[temp_w*0 +:temp_w];
assign v2119ibus[data_w*0 +:data_w] = c871obus[data_w*5 +:data_w];
assign c872ibus[temp_w*0 +:temp_w] = v486obus[temp_w*4 +:temp_w];
assign v486ibus[data_w*4 +:data_w] = c872obus[data_w*0 +:data_w];
assign c872ibus[temp_w*1 +:temp_w] = v739obus[temp_w*4 +:temp_w];
assign v739ibus[data_w*4 +:data_w] = c872obus[data_w*1 +:data_w];
assign c872ibus[temp_w*2 +:temp_w] = v1038obus[temp_w*2 +:temp_w];
assign v1038ibus[data_w*2 +:data_w] = c872obus[data_w*2 +:data_w];
assign c872ibus[temp_w*3 +:temp_w] = v1136obus[temp_w*4 +:temp_w];
assign v1136ibus[data_w*4 +:data_w] = c872obus[data_w*3 +:data_w];
assign c872ibus[temp_w*4 +:temp_w] = v2024obus[temp_w*1 +:temp_w];
assign v2024ibus[data_w*1 +:data_w] = c872obus[data_w*4 +:data_w];
assign c872ibus[temp_w*5 +:temp_w] = v2120obus[temp_w*0 +:temp_w];
assign v2120ibus[data_w*0 +:data_w] = c872obus[data_w*5 +:data_w];
assign c873ibus[temp_w*0 +:temp_w] = v487obus[temp_w*4 +:temp_w];
assign v487ibus[data_w*4 +:data_w] = c873obus[data_w*0 +:data_w];
assign c873ibus[temp_w*1 +:temp_w] = v740obus[temp_w*4 +:temp_w];
assign v740ibus[data_w*4 +:data_w] = c873obus[data_w*1 +:data_w];
assign c873ibus[temp_w*2 +:temp_w] = v1039obus[temp_w*2 +:temp_w];
assign v1039ibus[data_w*2 +:data_w] = c873obus[data_w*2 +:data_w];
assign c873ibus[temp_w*3 +:temp_w] = v1137obus[temp_w*4 +:temp_w];
assign v1137ibus[data_w*4 +:data_w] = c873obus[data_w*3 +:data_w];
assign c873ibus[temp_w*4 +:temp_w] = v2025obus[temp_w*1 +:temp_w];
assign v2025ibus[data_w*1 +:data_w] = c873obus[data_w*4 +:data_w];
assign c873ibus[temp_w*5 +:temp_w] = v2121obus[temp_w*0 +:temp_w];
assign v2121ibus[data_w*0 +:data_w] = c873obus[data_w*5 +:data_w];
assign c874ibus[temp_w*0 +:temp_w] = v488obus[temp_w*4 +:temp_w];
assign v488ibus[data_w*4 +:data_w] = c874obus[data_w*0 +:data_w];
assign c874ibus[temp_w*1 +:temp_w] = v741obus[temp_w*4 +:temp_w];
assign v741ibus[data_w*4 +:data_w] = c874obus[data_w*1 +:data_w];
assign c874ibus[temp_w*2 +:temp_w] = v1040obus[temp_w*2 +:temp_w];
assign v1040ibus[data_w*2 +:data_w] = c874obus[data_w*2 +:data_w];
assign c874ibus[temp_w*3 +:temp_w] = v1138obus[temp_w*4 +:temp_w];
assign v1138ibus[data_w*4 +:data_w] = c874obus[data_w*3 +:data_w];
assign c874ibus[temp_w*4 +:temp_w] = v2026obus[temp_w*1 +:temp_w];
assign v2026ibus[data_w*1 +:data_w] = c874obus[data_w*4 +:data_w];
assign c874ibus[temp_w*5 +:temp_w] = v2122obus[temp_w*0 +:temp_w];
assign v2122ibus[data_w*0 +:data_w] = c874obus[data_w*5 +:data_w];
assign c875ibus[temp_w*0 +:temp_w] = v489obus[temp_w*4 +:temp_w];
assign v489ibus[data_w*4 +:data_w] = c875obus[data_w*0 +:data_w];
assign c875ibus[temp_w*1 +:temp_w] = v742obus[temp_w*4 +:temp_w];
assign v742ibus[data_w*4 +:data_w] = c875obus[data_w*1 +:data_w];
assign c875ibus[temp_w*2 +:temp_w] = v1041obus[temp_w*2 +:temp_w];
assign v1041ibus[data_w*2 +:data_w] = c875obus[data_w*2 +:data_w];
assign c875ibus[temp_w*3 +:temp_w] = v1139obus[temp_w*4 +:temp_w];
assign v1139ibus[data_w*4 +:data_w] = c875obus[data_w*3 +:data_w];
assign c875ibus[temp_w*4 +:temp_w] = v2027obus[temp_w*1 +:temp_w];
assign v2027ibus[data_w*1 +:data_w] = c875obus[data_w*4 +:data_w];
assign c875ibus[temp_w*5 +:temp_w] = v2123obus[temp_w*0 +:temp_w];
assign v2123ibus[data_w*0 +:data_w] = c875obus[data_w*5 +:data_w];
assign c876ibus[temp_w*0 +:temp_w] = v490obus[temp_w*4 +:temp_w];
assign v490ibus[data_w*4 +:data_w] = c876obus[data_w*0 +:data_w];
assign c876ibus[temp_w*1 +:temp_w] = v743obus[temp_w*4 +:temp_w];
assign v743ibus[data_w*4 +:data_w] = c876obus[data_w*1 +:data_w];
assign c876ibus[temp_w*2 +:temp_w] = v1042obus[temp_w*2 +:temp_w];
assign v1042ibus[data_w*2 +:data_w] = c876obus[data_w*2 +:data_w];
assign c876ibus[temp_w*3 +:temp_w] = v1140obus[temp_w*4 +:temp_w];
assign v1140ibus[data_w*4 +:data_w] = c876obus[data_w*3 +:data_w];
assign c876ibus[temp_w*4 +:temp_w] = v2028obus[temp_w*1 +:temp_w];
assign v2028ibus[data_w*1 +:data_w] = c876obus[data_w*4 +:data_w];
assign c876ibus[temp_w*5 +:temp_w] = v2124obus[temp_w*0 +:temp_w];
assign v2124ibus[data_w*0 +:data_w] = c876obus[data_w*5 +:data_w];
assign c877ibus[temp_w*0 +:temp_w] = v491obus[temp_w*4 +:temp_w];
assign v491ibus[data_w*4 +:data_w] = c877obus[data_w*0 +:data_w];
assign c877ibus[temp_w*1 +:temp_w] = v744obus[temp_w*4 +:temp_w];
assign v744ibus[data_w*4 +:data_w] = c877obus[data_w*1 +:data_w];
assign c877ibus[temp_w*2 +:temp_w] = v1043obus[temp_w*2 +:temp_w];
assign v1043ibus[data_w*2 +:data_w] = c877obus[data_w*2 +:data_w];
assign c877ibus[temp_w*3 +:temp_w] = v1141obus[temp_w*4 +:temp_w];
assign v1141ibus[data_w*4 +:data_w] = c877obus[data_w*3 +:data_w];
assign c877ibus[temp_w*4 +:temp_w] = v2029obus[temp_w*1 +:temp_w];
assign v2029ibus[data_w*1 +:data_w] = c877obus[data_w*4 +:data_w];
assign c877ibus[temp_w*5 +:temp_w] = v2125obus[temp_w*0 +:temp_w];
assign v2125ibus[data_w*0 +:data_w] = c877obus[data_w*5 +:data_w];
assign c878ibus[temp_w*0 +:temp_w] = v492obus[temp_w*4 +:temp_w];
assign v492ibus[data_w*4 +:data_w] = c878obus[data_w*0 +:data_w];
assign c878ibus[temp_w*1 +:temp_w] = v745obus[temp_w*4 +:temp_w];
assign v745ibus[data_w*4 +:data_w] = c878obus[data_w*1 +:data_w];
assign c878ibus[temp_w*2 +:temp_w] = v1044obus[temp_w*2 +:temp_w];
assign v1044ibus[data_w*2 +:data_w] = c878obus[data_w*2 +:data_w];
assign c878ibus[temp_w*3 +:temp_w] = v1142obus[temp_w*4 +:temp_w];
assign v1142ibus[data_w*4 +:data_w] = c878obus[data_w*3 +:data_w];
assign c878ibus[temp_w*4 +:temp_w] = v2030obus[temp_w*1 +:temp_w];
assign v2030ibus[data_w*1 +:data_w] = c878obus[data_w*4 +:data_w];
assign c878ibus[temp_w*5 +:temp_w] = v2126obus[temp_w*0 +:temp_w];
assign v2126ibus[data_w*0 +:data_w] = c878obus[data_w*5 +:data_w];
assign c879ibus[temp_w*0 +:temp_w] = v493obus[temp_w*4 +:temp_w];
assign v493ibus[data_w*4 +:data_w] = c879obus[data_w*0 +:data_w];
assign c879ibus[temp_w*1 +:temp_w] = v746obus[temp_w*4 +:temp_w];
assign v746ibus[data_w*4 +:data_w] = c879obus[data_w*1 +:data_w];
assign c879ibus[temp_w*2 +:temp_w] = v1045obus[temp_w*2 +:temp_w];
assign v1045ibus[data_w*2 +:data_w] = c879obus[data_w*2 +:data_w];
assign c879ibus[temp_w*3 +:temp_w] = v1143obus[temp_w*4 +:temp_w];
assign v1143ibus[data_w*4 +:data_w] = c879obus[data_w*3 +:data_w];
assign c879ibus[temp_w*4 +:temp_w] = v2031obus[temp_w*1 +:temp_w];
assign v2031ibus[data_w*1 +:data_w] = c879obus[data_w*4 +:data_w];
assign c879ibus[temp_w*5 +:temp_w] = v2127obus[temp_w*0 +:temp_w];
assign v2127ibus[data_w*0 +:data_w] = c879obus[data_w*5 +:data_w];
assign c880ibus[temp_w*0 +:temp_w] = v494obus[temp_w*4 +:temp_w];
assign v494ibus[data_w*4 +:data_w] = c880obus[data_w*0 +:data_w];
assign c880ibus[temp_w*1 +:temp_w] = v747obus[temp_w*4 +:temp_w];
assign v747ibus[data_w*4 +:data_w] = c880obus[data_w*1 +:data_w];
assign c880ibus[temp_w*2 +:temp_w] = v1046obus[temp_w*2 +:temp_w];
assign v1046ibus[data_w*2 +:data_w] = c880obus[data_w*2 +:data_w];
assign c880ibus[temp_w*3 +:temp_w] = v1144obus[temp_w*4 +:temp_w];
assign v1144ibus[data_w*4 +:data_w] = c880obus[data_w*3 +:data_w];
assign c880ibus[temp_w*4 +:temp_w] = v2032obus[temp_w*1 +:temp_w];
assign v2032ibus[data_w*1 +:data_w] = c880obus[data_w*4 +:data_w];
assign c880ibus[temp_w*5 +:temp_w] = v2128obus[temp_w*0 +:temp_w];
assign v2128ibus[data_w*0 +:data_w] = c880obus[data_w*5 +:data_w];
assign c881ibus[temp_w*0 +:temp_w] = v495obus[temp_w*4 +:temp_w];
assign v495ibus[data_w*4 +:data_w] = c881obus[data_w*0 +:data_w];
assign c881ibus[temp_w*1 +:temp_w] = v748obus[temp_w*4 +:temp_w];
assign v748ibus[data_w*4 +:data_w] = c881obus[data_w*1 +:data_w];
assign c881ibus[temp_w*2 +:temp_w] = v1047obus[temp_w*2 +:temp_w];
assign v1047ibus[data_w*2 +:data_w] = c881obus[data_w*2 +:data_w];
assign c881ibus[temp_w*3 +:temp_w] = v1145obus[temp_w*4 +:temp_w];
assign v1145ibus[data_w*4 +:data_w] = c881obus[data_w*3 +:data_w];
assign c881ibus[temp_w*4 +:temp_w] = v2033obus[temp_w*1 +:temp_w];
assign v2033ibus[data_w*1 +:data_w] = c881obus[data_w*4 +:data_w];
assign c881ibus[temp_w*5 +:temp_w] = v2129obus[temp_w*0 +:temp_w];
assign v2129ibus[data_w*0 +:data_w] = c881obus[data_w*5 +:data_w];
assign c882ibus[temp_w*0 +:temp_w] = v496obus[temp_w*4 +:temp_w];
assign v496ibus[data_w*4 +:data_w] = c882obus[data_w*0 +:data_w];
assign c882ibus[temp_w*1 +:temp_w] = v749obus[temp_w*4 +:temp_w];
assign v749ibus[data_w*4 +:data_w] = c882obus[data_w*1 +:data_w];
assign c882ibus[temp_w*2 +:temp_w] = v1048obus[temp_w*2 +:temp_w];
assign v1048ibus[data_w*2 +:data_w] = c882obus[data_w*2 +:data_w];
assign c882ibus[temp_w*3 +:temp_w] = v1146obus[temp_w*4 +:temp_w];
assign v1146ibus[data_w*4 +:data_w] = c882obus[data_w*3 +:data_w];
assign c882ibus[temp_w*4 +:temp_w] = v2034obus[temp_w*1 +:temp_w];
assign v2034ibus[data_w*1 +:data_w] = c882obus[data_w*4 +:data_w];
assign c882ibus[temp_w*5 +:temp_w] = v2130obus[temp_w*0 +:temp_w];
assign v2130ibus[data_w*0 +:data_w] = c882obus[data_w*5 +:data_w];
assign c883ibus[temp_w*0 +:temp_w] = v497obus[temp_w*4 +:temp_w];
assign v497ibus[data_w*4 +:data_w] = c883obus[data_w*0 +:data_w];
assign c883ibus[temp_w*1 +:temp_w] = v750obus[temp_w*4 +:temp_w];
assign v750ibus[data_w*4 +:data_w] = c883obus[data_w*1 +:data_w];
assign c883ibus[temp_w*2 +:temp_w] = v1049obus[temp_w*2 +:temp_w];
assign v1049ibus[data_w*2 +:data_w] = c883obus[data_w*2 +:data_w];
assign c883ibus[temp_w*3 +:temp_w] = v1147obus[temp_w*4 +:temp_w];
assign v1147ibus[data_w*4 +:data_w] = c883obus[data_w*3 +:data_w];
assign c883ibus[temp_w*4 +:temp_w] = v2035obus[temp_w*1 +:temp_w];
assign v2035ibus[data_w*1 +:data_w] = c883obus[data_w*4 +:data_w];
assign c883ibus[temp_w*5 +:temp_w] = v2131obus[temp_w*0 +:temp_w];
assign v2131ibus[data_w*0 +:data_w] = c883obus[data_w*5 +:data_w];
assign c884ibus[temp_w*0 +:temp_w] = v498obus[temp_w*4 +:temp_w];
assign v498ibus[data_w*4 +:data_w] = c884obus[data_w*0 +:data_w];
assign c884ibus[temp_w*1 +:temp_w] = v751obus[temp_w*4 +:temp_w];
assign v751ibus[data_w*4 +:data_w] = c884obus[data_w*1 +:data_w];
assign c884ibus[temp_w*2 +:temp_w] = v1050obus[temp_w*2 +:temp_w];
assign v1050ibus[data_w*2 +:data_w] = c884obus[data_w*2 +:data_w];
assign c884ibus[temp_w*3 +:temp_w] = v1148obus[temp_w*4 +:temp_w];
assign v1148ibus[data_w*4 +:data_w] = c884obus[data_w*3 +:data_w];
assign c884ibus[temp_w*4 +:temp_w] = v2036obus[temp_w*1 +:temp_w];
assign v2036ibus[data_w*1 +:data_w] = c884obus[data_w*4 +:data_w];
assign c884ibus[temp_w*5 +:temp_w] = v2132obus[temp_w*0 +:temp_w];
assign v2132ibus[data_w*0 +:data_w] = c884obus[data_w*5 +:data_w];
assign c885ibus[temp_w*0 +:temp_w] = v499obus[temp_w*4 +:temp_w];
assign v499ibus[data_w*4 +:data_w] = c885obus[data_w*0 +:data_w];
assign c885ibus[temp_w*1 +:temp_w] = v752obus[temp_w*4 +:temp_w];
assign v752ibus[data_w*4 +:data_w] = c885obus[data_w*1 +:data_w];
assign c885ibus[temp_w*2 +:temp_w] = v1051obus[temp_w*2 +:temp_w];
assign v1051ibus[data_w*2 +:data_w] = c885obus[data_w*2 +:data_w];
assign c885ibus[temp_w*3 +:temp_w] = v1149obus[temp_w*4 +:temp_w];
assign v1149ibus[data_w*4 +:data_w] = c885obus[data_w*3 +:data_w];
assign c885ibus[temp_w*4 +:temp_w] = v2037obus[temp_w*1 +:temp_w];
assign v2037ibus[data_w*1 +:data_w] = c885obus[data_w*4 +:data_w];
assign c885ibus[temp_w*5 +:temp_w] = v2133obus[temp_w*0 +:temp_w];
assign v2133ibus[data_w*0 +:data_w] = c885obus[data_w*5 +:data_w];
assign c886ibus[temp_w*0 +:temp_w] = v500obus[temp_w*4 +:temp_w];
assign v500ibus[data_w*4 +:data_w] = c886obus[data_w*0 +:data_w];
assign c886ibus[temp_w*1 +:temp_w] = v753obus[temp_w*4 +:temp_w];
assign v753ibus[data_w*4 +:data_w] = c886obus[data_w*1 +:data_w];
assign c886ibus[temp_w*2 +:temp_w] = v1052obus[temp_w*2 +:temp_w];
assign v1052ibus[data_w*2 +:data_w] = c886obus[data_w*2 +:data_w];
assign c886ibus[temp_w*3 +:temp_w] = v1150obus[temp_w*4 +:temp_w];
assign v1150ibus[data_w*4 +:data_w] = c886obus[data_w*3 +:data_w];
assign c886ibus[temp_w*4 +:temp_w] = v2038obus[temp_w*1 +:temp_w];
assign v2038ibus[data_w*1 +:data_w] = c886obus[data_w*4 +:data_w];
assign c886ibus[temp_w*5 +:temp_w] = v2134obus[temp_w*0 +:temp_w];
assign v2134ibus[data_w*0 +:data_w] = c886obus[data_w*5 +:data_w];
assign c887ibus[temp_w*0 +:temp_w] = v501obus[temp_w*4 +:temp_w];
assign v501ibus[data_w*4 +:data_w] = c887obus[data_w*0 +:data_w];
assign c887ibus[temp_w*1 +:temp_w] = v754obus[temp_w*4 +:temp_w];
assign v754ibus[data_w*4 +:data_w] = c887obus[data_w*1 +:data_w];
assign c887ibus[temp_w*2 +:temp_w] = v1053obus[temp_w*2 +:temp_w];
assign v1053ibus[data_w*2 +:data_w] = c887obus[data_w*2 +:data_w];
assign c887ibus[temp_w*3 +:temp_w] = v1151obus[temp_w*4 +:temp_w];
assign v1151ibus[data_w*4 +:data_w] = c887obus[data_w*3 +:data_w];
assign c887ibus[temp_w*4 +:temp_w] = v2039obus[temp_w*1 +:temp_w];
assign v2039ibus[data_w*1 +:data_w] = c887obus[data_w*4 +:data_w];
assign c887ibus[temp_w*5 +:temp_w] = v2135obus[temp_w*0 +:temp_w];
assign v2135ibus[data_w*0 +:data_w] = c887obus[data_w*5 +:data_w];
assign c888ibus[temp_w*0 +:temp_w] = v502obus[temp_w*4 +:temp_w];
assign v502ibus[data_w*4 +:data_w] = c888obus[data_w*0 +:data_w];
assign c888ibus[temp_w*1 +:temp_w] = v755obus[temp_w*4 +:temp_w];
assign v755ibus[data_w*4 +:data_w] = c888obus[data_w*1 +:data_w];
assign c888ibus[temp_w*2 +:temp_w] = v1054obus[temp_w*2 +:temp_w];
assign v1054ibus[data_w*2 +:data_w] = c888obus[data_w*2 +:data_w];
assign c888ibus[temp_w*3 +:temp_w] = v1056obus[temp_w*4 +:temp_w];
assign v1056ibus[data_w*4 +:data_w] = c888obus[data_w*3 +:data_w];
assign c888ibus[temp_w*4 +:temp_w] = v2040obus[temp_w*1 +:temp_w];
assign v2040ibus[data_w*1 +:data_w] = c888obus[data_w*4 +:data_w];
assign c888ibus[temp_w*5 +:temp_w] = v2136obus[temp_w*0 +:temp_w];
assign v2136ibus[data_w*0 +:data_w] = c888obus[data_w*5 +:data_w];
assign c889ibus[temp_w*0 +:temp_w] = v503obus[temp_w*4 +:temp_w];
assign v503ibus[data_w*4 +:data_w] = c889obus[data_w*0 +:data_w];
assign c889ibus[temp_w*1 +:temp_w] = v756obus[temp_w*4 +:temp_w];
assign v756ibus[data_w*4 +:data_w] = c889obus[data_w*1 +:data_w];
assign c889ibus[temp_w*2 +:temp_w] = v1055obus[temp_w*2 +:temp_w];
assign v1055ibus[data_w*2 +:data_w] = c889obus[data_w*2 +:data_w];
assign c889ibus[temp_w*3 +:temp_w] = v1057obus[temp_w*4 +:temp_w];
assign v1057ibus[data_w*4 +:data_w] = c889obus[data_w*3 +:data_w];
assign c889ibus[temp_w*4 +:temp_w] = v2041obus[temp_w*1 +:temp_w];
assign v2041ibus[data_w*1 +:data_w] = c889obus[data_w*4 +:data_w];
assign c889ibus[temp_w*5 +:temp_w] = v2137obus[temp_w*0 +:temp_w];
assign v2137ibus[data_w*0 +:data_w] = c889obus[data_w*5 +:data_w];
assign c890ibus[temp_w*0 +:temp_w] = v504obus[temp_w*4 +:temp_w];
assign v504ibus[data_w*4 +:data_w] = c890obus[data_w*0 +:data_w];
assign c890ibus[temp_w*1 +:temp_w] = v757obus[temp_w*4 +:temp_w];
assign v757ibus[data_w*4 +:data_w] = c890obus[data_w*1 +:data_w];
assign c890ibus[temp_w*2 +:temp_w] = v960obus[temp_w*2 +:temp_w];
assign v960ibus[data_w*2 +:data_w] = c890obus[data_w*2 +:data_w];
assign c890ibus[temp_w*3 +:temp_w] = v1058obus[temp_w*4 +:temp_w];
assign v1058ibus[data_w*4 +:data_w] = c890obus[data_w*3 +:data_w];
assign c890ibus[temp_w*4 +:temp_w] = v2042obus[temp_w*1 +:temp_w];
assign v2042ibus[data_w*1 +:data_w] = c890obus[data_w*4 +:data_w];
assign c890ibus[temp_w*5 +:temp_w] = v2138obus[temp_w*0 +:temp_w];
assign v2138ibus[data_w*0 +:data_w] = c890obus[data_w*5 +:data_w];
assign c891ibus[temp_w*0 +:temp_w] = v505obus[temp_w*4 +:temp_w];
assign v505ibus[data_w*4 +:data_w] = c891obus[data_w*0 +:data_w];
assign c891ibus[temp_w*1 +:temp_w] = v758obus[temp_w*4 +:temp_w];
assign v758ibus[data_w*4 +:data_w] = c891obus[data_w*1 +:data_w];
assign c891ibus[temp_w*2 +:temp_w] = v961obus[temp_w*2 +:temp_w];
assign v961ibus[data_w*2 +:data_w] = c891obus[data_w*2 +:data_w];
assign c891ibus[temp_w*3 +:temp_w] = v1059obus[temp_w*4 +:temp_w];
assign v1059ibus[data_w*4 +:data_w] = c891obus[data_w*3 +:data_w];
assign c891ibus[temp_w*4 +:temp_w] = v2043obus[temp_w*1 +:temp_w];
assign v2043ibus[data_w*1 +:data_w] = c891obus[data_w*4 +:data_w];
assign c891ibus[temp_w*5 +:temp_w] = v2139obus[temp_w*0 +:temp_w];
assign v2139ibus[data_w*0 +:data_w] = c891obus[data_w*5 +:data_w];
assign c892ibus[temp_w*0 +:temp_w] = v506obus[temp_w*4 +:temp_w];
assign v506ibus[data_w*4 +:data_w] = c892obus[data_w*0 +:data_w];
assign c892ibus[temp_w*1 +:temp_w] = v759obus[temp_w*4 +:temp_w];
assign v759ibus[data_w*4 +:data_w] = c892obus[data_w*1 +:data_w];
assign c892ibus[temp_w*2 +:temp_w] = v962obus[temp_w*2 +:temp_w];
assign v962ibus[data_w*2 +:data_w] = c892obus[data_w*2 +:data_w];
assign c892ibus[temp_w*3 +:temp_w] = v1060obus[temp_w*4 +:temp_w];
assign v1060ibus[data_w*4 +:data_w] = c892obus[data_w*3 +:data_w];
assign c892ibus[temp_w*4 +:temp_w] = v2044obus[temp_w*1 +:temp_w];
assign v2044ibus[data_w*1 +:data_w] = c892obus[data_w*4 +:data_w];
assign c892ibus[temp_w*5 +:temp_w] = v2140obus[temp_w*0 +:temp_w];
assign v2140ibus[data_w*0 +:data_w] = c892obus[data_w*5 +:data_w];
assign c893ibus[temp_w*0 +:temp_w] = v507obus[temp_w*4 +:temp_w];
assign v507ibus[data_w*4 +:data_w] = c893obus[data_w*0 +:data_w];
assign c893ibus[temp_w*1 +:temp_w] = v760obus[temp_w*4 +:temp_w];
assign v760ibus[data_w*4 +:data_w] = c893obus[data_w*1 +:data_w];
assign c893ibus[temp_w*2 +:temp_w] = v963obus[temp_w*2 +:temp_w];
assign v963ibus[data_w*2 +:data_w] = c893obus[data_w*2 +:data_w];
assign c893ibus[temp_w*3 +:temp_w] = v1061obus[temp_w*4 +:temp_w];
assign v1061ibus[data_w*4 +:data_w] = c893obus[data_w*3 +:data_w];
assign c893ibus[temp_w*4 +:temp_w] = v2045obus[temp_w*1 +:temp_w];
assign v2045ibus[data_w*1 +:data_w] = c893obus[data_w*4 +:data_w];
assign c893ibus[temp_w*5 +:temp_w] = v2141obus[temp_w*0 +:temp_w];
assign v2141ibus[data_w*0 +:data_w] = c893obus[data_w*5 +:data_w];
assign c894ibus[temp_w*0 +:temp_w] = v508obus[temp_w*4 +:temp_w];
assign v508ibus[data_w*4 +:data_w] = c894obus[data_w*0 +:data_w];
assign c894ibus[temp_w*1 +:temp_w] = v761obus[temp_w*4 +:temp_w];
assign v761ibus[data_w*4 +:data_w] = c894obus[data_w*1 +:data_w];
assign c894ibus[temp_w*2 +:temp_w] = v964obus[temp_w*2 +:temp_w];
assign v964ibus[data_w*2 +:data_w] = c894obus[data_w*2 +:data_w];
assign c894ibus[temp_w*3 +:temp_w] = v1062obus[temp_w*4 +:temp_w];
assign v1062ibus[data_w*4 +:data_w] = c894obus[data_w*3 +:data_w];
assign c894ibus[temp_w*4 +:temp_w] = v2046obus[temp_w*1 +:temp_w];
assign v2046ibus[data_w*1 +:data_w] = c894obus[data_w*4 +:data_w];
assign c894ibus[temp_w*5 +:temp_w] = v2142obus[temp_w*0 +:temp_w];
assign v2142ibus[data_w*0 +:data_w] = c894obus[data_w*5 +:data_w];
assign c895ibus[temp_w*0 +:temp_w] = v509obus[temp_w*4 +:temp_w];
assign v509ibus[data_w*4 +:data_w] = c895obus[data_w*0 +:data_w];
assign c895ibus[temp_w*1 +:temp_w] = v762obus[temp_w*4 +:temp_w];
assign v762ibus[data_w*4 +:data_w] = c895obus[data_w*1 +:data_w];
assign c895ibus[temp_w*2 +:temp_w] = v965obus[temp_w*2 +:temp_w];
assign v965ibus[data_w*2 +:data_w] = c895obus[data_w*2 +:data_w];
assign c895ibus[temp_w*3 +:temp_w] = v1063obus[temp_w*4 +:temp_w];
assign v1063ibus[data_w*4 +:data_w] = c895obus[data_w*3 +:data_w];
assign c895ibus[temp_w*4 +:temp_w] = v2047obus[temp_w*1 +:temp_w];
assign v2047ibus[data_w*1 +:data_w] = c895obus[data_w*4 +:data_w];
assign c895ibus[temp_w*5 +:temp_w] = v2143obus[temp_w*0 +:temp_w];
assign v2143ibus[data_w*0 +:data_w] = c895obus[data_w*5 +:data_w];
assign c896ibus[temp_w*0 +:temp_w] = v510obus[temp_w*4 +:temp_w];
assign v510ibus[data_w*4 +:data_w] = c896obus[data_w*0 +:data_w];
assign c896ibus[temp_w*1 +:temp_w] = v763obus[temp_w*4 +:temp_w];
assign v763ibus[data_w*4 +:data_w] = c896obus[data_w*1 +:data_w];
assign c896ibus[temp_w*2 +:temp_w] = v966obus[temp_w*2 +:temp_w];
assign v966ibus[data_w*2 +:data_w] = c896obus[data_w*2 +:data_w];
assign c896ibus[temp_w*3 +:temp_w] = v1064obus[temp_w*4 +:temp_w];
assign v1064ibus[data_w*4 +:data_w] = c896obus[data_w*3 +:data_w];
assign c896ibus[temp_w*4 +:temp_w] = v2048obus[temp_w*1 +:temp_w];
assign v2048ibus[data_w*1 +:data_w] = c896obus[data_w*4 +:data_w];
assign c896ibus[temp_w*5 +:temp_w] = v2144obus[temp_w*0 +:temp_w];
assign v2144ibus[data_w*0 +:data_w] = c896obus[data_w*5 +:data_w];
assign c897ibus[temp_w*0 +:temp_w] = v511obus[temp_w*4 +:temp_w];
assign v511ibus[data_w*4 +:data_w] = c897obus[data_w*0 +:data_w];
assign c897ibus[temp_w*1 +:temp_w] = v764obus[temp_w*4 +:temp_w];
assign v764ibus[data_w*4 +:data_w] = c897obus[data_w*1 +:data_w];
assign c897ibus[temp_w*2 +:temp_w] = v967obus[temp_w*2 +:temp_w];
assign v967ibus[data_w*2 +:data_w] = c897obus[data_w*2 +:data_w];
assign c897ibus[temp_w*3 +:temp_w] = v1065obus[temp_w*4 +:temp_w];
assign v1065ibus[data_w*4 +:data_w] = c897obus[data_w*3 +:data_w];
assign c897ibus[temp_w*4 +:temp_w] = v2049obus[temp_w*1 +:temp_w];
assign v2049ibus[data_w*1 +:data_w] = c897obus[data_w*4 +:data_w];
assign c897ibus[temp_w*5 +:temp_w] = v2145obus[temp_w*0 +:temp_w];
assign v2145ibus[data_w*0 +:data_w] = c897obus[data_w*5 +:data_w];
assign c898ibus[temp_w*0 +:temp_w] = v512obus[temp_w*4 +:temp_w];
assign v512ibus[data_w*4 +:data_w] = c898obus[data_w*0 +:data_w];
assign c898ibus[temp_w*1 +:temp_w] = v765obus[temp_w*4 +:temp_w];
assign v765ibus[data_w*4 +:data_w] = c898obus[data_w*1 +:data_w];
assign c898ibus[temp_w*2 +:temp_w] = v968obus[temp_w*2 +:temp_w];
assign v968ibus[data_w*2 +:data_w] = c898obus[data_w*2 +:data_w];
assign c898ibus[temp_w*3 +:temp_w] = v1066obus[temp_w*4 +:temp_w];
assign v1066ibus[data_w*4 +:data_w] = c898obus[data_w*3 +:data_w];
assign c898ibus[temp_w*4 +:temp_w] = v2050obus[temp_w*1 +:temp_w];
assign v2050ibus[data_w*1 +:data_w] = c898obus[data_w*4 +:data_w];
assign c898ibus[temp_w*5 +:temp_w] = v2146obus[temp_w*0 +:temp_w];
assign v2146ibus[data_w*0 +:data_w] = c898obus[data_w*5 +:data_w];
assign c899ibus[temp_w*0 +:temp_w] = v513obus[temp_w*4 +:temp_w];
assign v513ibus[data_w*4 +:data_w] = c899obus[data_w*0 +:data_w];
assign c899ibus[temp_w*1 +:temp_w] = v766obus[temp_w*4 +:temp_w];
assign v766ibus[data_w*4 +:data_w] = c899obus[data_w*1 +:data_w];
assign c899ibus[temp_w*2 +:temp_w] = v969obus[temp_w*2 +:temp_w];
assign v969ibus[data_w*2 +:data_w] = c899obus[data_w*2 +:data_w];
assign c899ibus[temp_w*3 +:temp_w] = v1067obus[temp_w*4 +:temp_w];
assign v1067ibus[data_w*4 +:data_w] = c899obus[data_w*3 +:data_w];
assign c899ibus[temp_w*4 +:temp_w] = v2051obus[temp_w*1 +:temp_w];
assign v2051ibus[data_w*1 +:data_w] = c899obus[data_w*4 +:data_w];
assign c899ibus[temp_w*5 +:temp_w] = v2147obus[temp_w*0 +:temp_w];
assign v2147ibus[data_w*0 +:data_w] = c899obus[data_w*5 +:data_w];
assign c900ibus[temp_w*0 +:temp_w] = v514obus[temp_w*4 +:temp_w];
assign v514ibus[data_w*4 +:data_w] = c900obus[data_w*0 +:data_w];
assign c900ibus[temp_w*1 +:temp_w] = v767obus[temp_w*4 +:temp_w];
assign v767ibus[data_w*4 +:data_w] = c900obus[data_w*1 +:data_w];
assign c900ibus[temp_w*2 +:temp_w] = v970obus[temp_w*2 +:temp_w];
assign v970ibus[data_w*2 +:data_w] = c900obus[data_w*2 +:data_w];
assign c900ibus[temp_w*3 +:temp_w] = v1068obus[temp_w*4 +:temp_w];
assign v1068ibus[data_w*4 +:data_w] = c900obus[data_w*3 +:data_w];
assign c900ibus[temp_w*4 +:temp_w] = v2052obus[temp_w*1 +:temp_w];
assign v2052ibus[data_w*1 +:data_w] = c900obus[data_w*4 +:data_w];
assign c900ibus[temp_w*5 +:temp_w] = v2148obus[temp_w*0 +:temp_w];
assign v2148ibus[data_w*0 +:data_w] = c900obus[data_w*5 +:data_w];
assign c901ibus[temp_w*0 +:temp_w] = v515obus[temp_w*4 +:temp_w];
assign v515ibus[data_w*4 +:data_w] = c901obus[data_w*0 +:data_w];
assign c901ibus[temp_w*1 +:temp_w] = v672obus[temp_w*4 +:temp_w];
assign v672ibus[data_w*4 +:data_w] = c901obus[data_w*1 +:data_w];
assign c901ibus[temp_w*2 +:temp_w] = v971obus[temp_w*2 +:temp_w];
assign v971ibus[data_w*2 +:data_w] = c901obus[data_w*2 +:data_w];
assign c901ibus[temp_w*3 +:temp_w] = v1069obus[temp_w*4 +:temp_w];
assign v1069ibus[data_w*4 +:data_w] = c901obus[data_w*3 +:data_w];
assign c901ibus[temp_w*4 +:temp_w] = v2053obus[temp_w*1 +:temp_w];
assign v2053ibus[data_w*1 +:data_w] = c901obus[data_w*4 +:data_w];
assign c901ibus[temp_w*5 +:temp_w] = v2149obus[temp_w*0 +:temp_w];
assign v2149ibus[data_w*0 +:data_w] = c901obus[data_w*5 +:data_w];
assign c902ibus[temp_w*0 +:temp_w] = v516obus[temp_w*4 +:temp_w];
assign v516ibus[data_w*4 +:data_w] = c902obus[data_w*0 +:data_w];
assign c902ibus[temp_w*1 +:temp_w] = v673obus[temp_w*4 +:temp_w];
assign v673ibus[data_w*4 +:data_w] = c902obus[data_w*1 +:data_w];
assign c902ibus[temp_w*2 +:temp_w] = v972obus[temp_w*2 +:temp_w];
assign v972ibus[data_w*2 +:data_w] = c902obus[data_w*2 +:data_w];
assign c902ibus[temp_w*3 +:temp_w] = v1070obus[temp_w*4 +:temp_w];
assign v1070ibus[data_w*4 +:data_w] = c902obus[data_w*3 +:data_w];
assign c902ibus[temp_w*4 +:temp_w] = v2054obus[temp_w*1 +:temp_w];
assign v2054ibus[data_w*1 +:data_w] = c902obus[data_w*4 +:data_w];
assign c902ibus[temp_w*5 +:temp_w] = v2150obus[temp_w*0 +:temp_w];
assign v2150ibus[data_w*0 +:data_w] = c902obus[data_w*5 +:data_w];
assign c903ibus[temp_w*0 +:temp_w] = v517obus[temp_w*4 +:temp_w];
assign v517ibus[data_w*4 +:data_w] = c903obus[data_w*0 +:data_w];
assign c903ibus[temp_w*1 +:temp_w] = v674obus[temp_w*4 +:temp_w];
assign v674ibus[data_w*4 +:data_w] = c903obus[data_w*1 +:data_w];
assign c903ibus[temp_w*2 +:temp_w] = v973obus[temp_w*2 +:temp_w];
assign v973ibus[data_w*2 +:data_w] = c903obus[data_w*2 +:data_w];
assign c903ibus[temp_w*3 +:temp_w] = v1071obus[temp_w*4 +:temp_w];
assign v1071ibus[data_w*4 +:data_w] = c903obus[data_w*3 +:data_w];
assign c903ibus[temp_w*4 +:temp_w] = v2055obus[temp_w*1 +:temp_w];
assign v2055ibus[data_w*1 +:data_w] = c903obus[data_w*4 +:data_w];
assign c903ibus[temp_w*5 +:temp_w] = v2151obus[temp_w*0 +:temp_w];
assign v2151ibus[data_w*0 +:data_w] = c903obus[data_w*5 +:data_w];
assign c904ibus[temp_w*0 +:temp_w] = v518obus[temp_w*4 +:temp_w];
assign v518ibus[data_w*4 +:data_w] = c904obus[data_w*0 +:data_w];
assign c904ibus[temp_w*1 +:temp_w] = v675obus[temp_w*4 +:temp_w];
assign v675ibus[data_w*4 +:data_w] = c904obus[data_w*1 +:data_w];
assign c904ibus[temp_w*2 +:temp_w] = v974obus[temp_w*2 +:temp_w];
assign v974ibus[data_w*2 +:data_w] = c904obus[data_w*2 +:data_w];
assign c904ibus[temp_w*3 +:temp_w] = v1072obus[temp_w*4 +:temp_w];
assign v1072ibus[data_w*4 +:data_w] = c904obus[data_w*3 +:data_w];
assign c904ibus[temp_w*4 +:temp_w] = v2056obus[temp_w*1 +:temp_w];
assign v2056ibus[data_w*1 +:data_w] = c904obus[data_w*4 +:data_w];
assign c904ibus[temp_w*5 +:temp_w] = v2152obus[temp_w*0 +:temp_w];
assign v2152ibus[data_w*0 +:data_w] = c904obus[data_w*5 +:data_w];
assign c905ibus[temp_w*0 +:temp_w] = v519obus[temp_w*4 +:temp_w];
assign v519ibus[data_w*4 +:data_w] = c905obus[data_w*0 +:data_w];
assign c905ibus[temp_w*1 +:temp_w] = v676obus[temp_w*4 +:temp_w];
assign v676ibus[data_w*4 +:data_w] = c905obus[data_w*1 +:data_w];
assign c905ibus[temp_w*2 +:temp_w] = v975obus[temp_w*2 +:temp_w];
assign v975ibus[data_w*2 +:data_w] = c905obus[data_w*2 +:data_w];
assign c905ibus[temp_w*3 +:temp_w] = v1073obus[temp_w*4 +:temp_w];
assign v1073ibus[data_w*4 +:data_w] = c905obus[data_w*3 +:data_w];
assign c905ibus[temp_w*4 +:temp_w] = v2057obus[temp_w*1 +:temp_w];
assign v2057ibus[data_w*1 +:data_w] = c905obus[data_w*4 +:data_w];
assign c905ibus[temp_w*5 +:temp_w] = v2153obus[temp_w*0 +:temp_w];
assign v2153ibus[data_w*0 +:data_w] = c905obus[data_w*5 +:data_w];
assign c906ibus[temp_w*0 +:temp_w] = v520obus[temp_w*4 +:temp_w];
assign v520ibus[data_w*4 +:data_w] = c906obus[data_w*0 +:data_w];
assign c906ibus[temp_w*1 +:temp_w] = v677obus[temp_w*4 +:temp_w];
assign v677ibus[data_w*4 +:data_w] = c906obus[data_w*1 +:data_w];
assign c906ibus[temp_w*2 +:temp_w] = v976obus[temp_w*2 +:temp_w];
assign v976ibus[data_w*2 +:data_w] = c906obus[data_w*2 +:data_w];
assign c906ibus[temp_w*3 +:temp_w] = v1074obus[temp_w*4 +:temp_w];
assign v1074ibus[data_w*4 +:data_w] = c906obus[data_w*3 +:data_w];
assign c906ibus[temp_w*4 +:temp_w] = v2058obus[temp_w*1 +:temp_w];
assign v2058ibus[data_w*1 +:data_w] = c906obus[data_w*4 +:data_w];
assign c906ibus[temp_w*5 +:temp_w] = v2154obus[temp_w*0 +:temp_w];
assign v2154ibus[data_w*0 +:data_w] = c906obus[data_w*5 +:data_w];
assign c907ibus[temp_w*0 +:temp_w] = v521obus[temp_w*4 +:temp_w];
assign v521ibus[data_w*4 +:data_w] = c907obus[data_w*0 +:data_w];
assign c907ibus[temp_w*1 +:temp_w] = v678obus[temp_w*4 +:temp_w];
assign v678ibus[data_w*4 +:data_w] = c907obus[data_w*1 +:data_w];
assign c907ibus[temp_w*2 +:temp_w] = v977obus[temp_w*2 +:temp_w];
assign v977ibus[data_w*2 +:data_w] = c907obus[data_w*2 +:data_w];
assign c907ibus[temp_w*3 +:temp_w] = v1075obus[temp_w*4 +:temp_w];
assign v1075ibus[data_w*4 +:data_w] = c907obus[data_w*3 +:data_w];
assign c907ibus[temp_w*4 +:temp_w] = v2059obus[temp_w*1 +:temp_w];
assign v2059ibus[data_w*1 +:data_w] = c907obus[data_w*4 +:data_w];
assign c907ibus[temp_w*5 +:temp_w] = v2155obus[temp_w*0 +:temp_w];
assign v2155ibus[data_w*0 +:data_w] = c907obus[data_w*5 +:data_w];
assign c908ibus[temp_w*0 +:temp_w] = v522obus[temp_w*4 +:temp_w];
assign v522ibus[data_w*4 +:data_w] = c908obus[data_w*0 +:data_w];
assign c908ibus[temp_w*1 +:temp_w] = v679obus[temp_w*4 +:temp_w];
assign v679ibus[data_w*4 +:data_w] = c908obus[data_w*1 +:data_w];
assign c908ibus[temp_w*2 +:temp_w] = v978obus[temp_w*2 +:temp_w];
assign v978ibus[data_w*2 +:data_w] = c908obus[data_w*2 +:data_w];
assign c908ibus[temp_w*3 +:temp_w] = v1076obus[temp_w*4 +:temp_w];
assign v1076ibus[data_w*4 +:data_w] = c908obus[data_w*3 +:data_w];
assign c908ibus[temp_w*4 +:temp_w] = v2060obus[temp_w*1 +:temp_w];
assign v2060ibus[data_w*1 +:data_w] = c908obus[data_w*4 +:data_w];
assign c908ibus[temp_w*5 +:temp_w] = v2156obus[temp_w*0 +:temp_w];
assign v2156ibus[data_w*0 +:data_w] = c908obus[data_w*5 +:data_w];
assign c909ibus[temp_w*0 +:temp_w] = v523obus[temp_w*4 +:temp_w];
assign v523ibus[data_w*4 +:data_w] = c909obus[data_w*0 +:data_w];
assign c909ibus[temp_w*1 +:temp_w] = v680obus[temp_w*4 +:temp_w];
assign v680ibus[data_w*4 +:data_w] = c909obus[data_w*1 +:data_w];
assign c909ibus[temp_w*2 +:temp_w] = v979obus[temp_w*2 +:temp_w];
assign v979ibus[data_w*2 +:data_w] = c909obus[data_w*2 +:data_w];
assign c909ibus[temp_w*3 +:temp_w] = v1077obus[temp_w*4 +:temp_w];
assign v1077ibus[data_w*4 +:data_w] = c909obus[data_w*3 +:data_w];
assign c909ibus[temp_w*4 +:temp_w] = v2061obus[temp_w*1 +:temp_w];
assign v2061ibus[data_w*1 +:data_w] = c909obus[data_w*4 +:data_w];
assign c909ibus[temp_w*5 +:temp_w] = v2157obus[temp_w*0 +:temp_w];
assign v2157ibus[data_w*0 +:data_w] = c909obus[data_w*5 +:data_w];
assign c910ibus[temp_w*0 +:temp_w] = v524obus[temp_w*4 +:temp_w];
assign v524ibus[data_w*4 +:data_w] = c910obus[data_w*0 +:data_w];
assign c910ibus[temp_w*1 +:temp_w] = v681obus[temp_w*4 +:temp_w];
assign v681ibus[data_w*4 +:data_w] = c910obus[data_w*1 +:data_w];
assign c910ibus[temp_w*2 +:temp_w] = v980obus[temp_w*2 +:temp_w];
assign v980ibus[data_w*2 +:data_w] = c910obus[data_w*2 +:data_w];
assign c910ibus[temp_w*3 +:temp_w] = v1078obus[temp_w*4 +:temp_w];
assign v1078ibus[data_w*4 +:data_w] = c910obus[data_w*3 +:data_w];
assign c910ibus[temp_w*4 +:temp_w] = v2062obus[temp_w*1 +:temp_w];
assign v2062ibus[data_w*1 +:data_w] = c910obus[data_w*4 +:data_w];
assign c910ibus[temp_w*5 +:temp_w] = v2158obus[temp_w*0 +:temp_w];
assign v2158ibus[data_w*0 +:data_w] = c910obus[data_w*5 +:data_w];
assign c911ibus[temp_w*0 +:temp_w] = v525obus[temp_w*4 +:temp_w];
assign v525ibus[data_w*4 +:data_w] = c911obus[data_w*0 +:data_w];
assign c911ibus[temp_w*1 +:temp_w] = v682obus[temp_w*4 +:temp_w];
assign v682ibus[data_w*4 +:data_w] = c911obus[data_w*1 +:data_w];
assign c911ibus[temp_w*2 +:temp_w] = v981obus[temp_w*2 +:temp_w];
assign v981ibus[data_w*2 +:data_w] = c911obus[data_w*2 +:data_w];
assign c911ibus[temp_w*3 +:temp_w] = v1079obus[temp_w*4 +:temp_w];
assign v1079ibus[data_w*4 +:data_w] = c911obus[data_w*3 +:data_w];
assign c911ibus[temp_w*4 +:temp_w] = v2063obus[temp_w*1 +:temp_w];
assign v2063ibus[data_w*1 +:data_w] = c911obus[data_w*4 +:data_w];
assign c911ibus[temp_w*5 +:temp_w] = v2159obus[temp_w*0 +:temp_w];
assign v2159ibus[data_w*0 +:data_w] = c911obus[data_w*5 +:data_w];
assign c912ibus[temp_w*0 +:temp_w] = v526obus[temp_w*4 +:temp_w];
assign v526ibus[data_w*4 +:data_w] = c912obus[data_w*0 +:data_w];
assign c912ibus[temp_w*1 +:temp_w] = v683obus[temp_w*4 +:temp_w];
assign v683ibus[data_w*4 +:data_w] = c912obus[data_w*1 +:data_w];
assign c912ibus[temp_w*2 +:temp_w] = v982obus[temp_w*2 +:temp_w];
assign v982ibus[data_w*2 +:data_w] = c912obus[data_w*2 +:data_w];
assign c912ibus[temp_w*3 +:temp_w] = v1080obus[temp_w*4 +:temp_w];
assign v1080ibus[data_w*4 +:data_w] = c912obus[data_w*3 +:data_w];
assign c912ibus[temp_w*4 +:temp_w] = v2064obus[temp_w*1 +:temp_w];
assign v2064ibus[data_w*1 +:data_w] = c912obus[data_w*4 +:data_w];
assign c912ibus[temp_w*5 +:temp_w] = v2160obus[temp_w*0 +:temp_w];
assign v2160ibus[data_w*0 +:data_w] = c912obus[data_w*5 +:data_w];
assign c913ibus[temp_w*0 +:temp_w] = v527obus[temp_w*4 +:temp_w];
assign v527ibus[data_w*4 +:data_w] = c913obus[data_w*0 +:data_w];
assign c913ibus[temp_w*1 +:temp_w] = v684obus[temp_w*4 +:temp_w];
assign v684ibus[data_w*4 +:data_w] = c913obus[data_w*1 +:data_w];
assign c913ibus[temp_w*2 +:temp_w] = v983obus[temp_w*2 +:temp_w];
assign v983ibus[data_w*2 +:data_w] = c913obus[data_w*2 +:data_w];
assign c913ibus[temp_w*3 +:temp_w] = v1081obus[temp_w*4 +:temp_w];
assign v1081ibus[data_w*4 +:data_w] = c913obus[data_w*3 +:data_w];
assign c913ibus[temp_w*4 +:temp_w] = v2065obus[temp_w*1 +:temp_w];
assign v2065ibus[data_w*1 +:data_w] = c913obus[data_w*4 +:data_w];
assign c913ibus[temp_w*5 +:temp_w] = v2161obus[temp_w*0 +:temp_w];
assign v2161ibus[data_w*0 +:data_w] = c913obus[data_w*5 +:data_w];
assign c914ibus[temp_w*0 +:temp_w] = v528obus[temp_w*4 +:temp_w];
assign v528ibus[data_w*4 +:data_w] = c914obus[data_w*0 +:data_w];
assign c914ibus[temp_w*1 +:temp_w] = v685obus[temp_w*4 +:temp_w];
assign v685ibus[data_w*4 +:data_w] = c914obus[data_w*1 +:data_w];
assign c914ibus[temp_w*2 +:temp_w] = v984obus[temp_w*2 +:temp_w];
assign v984ibus[data_w*2 +:data_w] = c914obus[data_w*2 +:data_w];
assign c914ibus[temp_w*3 +:temp_w] = v1082obus[temp_w*4 +:temp_w];
assign v1082ibus[data_w*4 +:data_w] = c914obus[data_w*3 +:data_w];
assign c914ibus[temp_w*4 +:temp_w] = v2066obus[temp_w*1 +:temp_w];
assign v2066ibus[data_w*1 +:data_w] = c914obus[data_w*4 +:data_w];
assign c914ibus[temp_w*5 +:temp_w] = v2162obus[temp_w*0 +:temp_w];
assign v2162ibus[data_w*0 +:data_w] = c914obus[data_w*5 +:data_w];
assign c915ibus[temp_w*0 +:temp_w] = v529obus[temp_w*4 +:temp_w];
assign v529ibus[data_w*4 +:data_w] = c915obus[data_w*0 +:data_w];
assign c915ibus[temp_w*1 +:temp_w] = v686obus[temp_w*4 +:temp_w];
assign v686ibus[data_w*4 +:data_w] = c915obus[data_w*1 +:data_w];
assign c915ibus[temp_w*2 +:temp_w] = v985obus[temp_w*2 +:temp_w];
assign v985ibus[data_w*2 +:data_w] = c915obus[data_w*2 +:data_w];
assign c915ibus[temp_w*3 +:temp_w] = v1083obus[temp_w*4 +:temp_w];
assign v1083ibus[data_w*4 +:data_w] = c915obus[data_w*3 +:data_w];
assign c915ibus[temp_w*4 +:temp_w] = v2067obus[temp_w*1 +:temp_w];
assign v2067ibus[data_w*1 +:data_w] = c915obus[data_w*4 +:data_w];
assign c915ibus[temp_w*5 +:temp_w] = v2163obus[temp_w*0 +:temp_w];
assign v2163ibus[data_w*0 +:data_w] = c915obus[data_w*5 +:data_w];
assign c916ibus[temp_w*0 +:temp_w] = v530obus[temp_w*4 +:temp_w];
assign v530ibus[data_w*4 +:data_w] = c916obus[data_w*0 +:data_w];
assign c916ibus[temp_w*1 +:temp_w] = v687obus[temp_w*4 +:temp_w];
assign v687ibus[data_w*4 +:data_w] = c916obus[data_w*1 +:data_w];
assign c916ibus[temp_w*2 +:temp_w] = v986obus[temp_w*2 +:temp_w];
assign v986ibus[data_w*2 +:data_w] = c916obus[data_w*2 +:data_w];
assign c916ibus[temp_w*3 +:temp_w] = v1084obus[temp_w*4 +:temp_w];
assign v1084ibus[data_w*4 +:data_w] = c916obus[data_w*3 +:data_w];
assign c916ibus[temp_w*4 +:temp_w] = v2068obus[temp_w*1 +:temp_w];
assign v2068ibus[data_w*1 +:data_w] = c916obus[data_w*4 +:data_w];
assign c916ibus[temp_w*5 +:temp_w] = v2164obus[temp_w*0 +:temp_w];
assign v2164ibus[data_w*0 +:data_w] = c916obus[data_w*5 +:data_w];
assign c917ibus[temp_w*0 +:temp_w] = v531obus[temp_w*4 +:temp_w];
assign v531ibus[data_w*4 +:data_w] = c917obus[data_w*0 +:data_w];
assign c917ibus[temp_w*1 +:temp_w] = v688obus[temp_w*4 +:temp_w];
assign v688ibus[data_w*4 +:data_w] = c917obus[data_w*1 +:data_w];
assign c917ibus[temp_w*2 +:temp_w] = v987obus[temp_w*2 +:temp_w];
assign v987ibus[data_w*2 +:data_w] = c917obus[data_w*2 +:data_w];
assign c917ibus[temp_w*3 +:temp_w] = v1085obus[temp_w*4 +:temp_w];
assign v1085ibus[data_w*4 +:data_w] = c917obus[data_w*3 +:data_w];
assign c917ibus[temp_w*4 +:temp_w] = v2069obus[temp_w*1 +:temp_w];
assign v2069ibus[data_w*1 +:data_w] = c917obus[data_w*4 +:data_w];
assign c917ibus[temp_w*5 +:temp_w] = v2165obus[temp_w*0 +:temp_w];
assign v2165ibus[data_w*0 +:data_w] = c917obus[data_w*5 +:data_w];
assign c918ibus[temp_w*0 +:temp_w] = v532obus[temp_w*4 +:temp_w];
assign v532ibus[data_w*4 +:data_w] = c918obus[data_w*0 +:data_w];
assign c918ibus[temp_w*1 +:temp_w] = v689obus[temp_w*4 +:temp_w];
assign v689ibus[data_w*4 +:data_w] = c918obus[data_w*1 +:data_w];
assign c918ibus[temp_w*2 +:temp_w] = v988obus[temp_w*2 +:temp_w];
assign v988ibus[data_w*2 +:data_w] = c918obus[data_w*2 +:data_w];
assign c918ibus[temp_w*3 +:temp_w] = v1086obus[temp_w*4 +:temp_w];
assign v1086ibus[data_w*4 +:data_w] = c918obus[data_w*3 +:data_w];
assign c918ibus[temp_w*4 +:temp_w] = v2070obus[temp_w*1 +:temp_w];
assign v2070ibus[data_w*1 +:data_w] = c918obus[data_w*4 +:data_w];
assign c918ibus[temp_w*5 +:temp_w] = v2166obus[temp_w*0 +:temp_w];
assign v2166ibus[data_w*0 +:data_w] = c918obus[data_w*5 +:data_w];
assign c919ibus[temp_w*0 +:temp_w] = v533obus[temp_w*4 +:temp_w];
assign v533ibus[data_w*4 +:data_w] = c919obus[data_w*0 +:data_w];
assign c919ibus[temp_w*1 +:temp_w] = v690obus[temp_w*4 +:temp_w];
assign v690ibus[data_w*4 +:data_w] = c919obus[data_w*1 +:data_w];
assign c919ibus[temp_w*2 +:temp_w] = v989obus[temp_w*2 +:temp_w];
assign v989ibus[data_w*2 +:data_w] = c919obus[data_w*2 +:data_w];
assign c919ibus[temp_w*3 +:temp_w] = v1087obus[temp_w*4 +:temp_w];
assign v1087ibus[data_w*4 +:data_w] = c919obus[data_w*3 +:data_w];
assign c919ibus[temp_w*4 +:temp_w] = v2071obus[temp_w*1 +:temp_w];
assign v2071ibus[data_w*1 +:data_w] = c919obus[data_w*4 +:data_w];
assign c919ibus[temp_w*5 +:temp_w] = v2167obus[temp_w*0 +:temp_w];
assign v2167ibus[data_w*0 +:data_w] = c919obus[data_w*5 +:data_w];
assign c920ibus[temp_w*0 +:temp_w] = v534obus[temp_w*4 +:temp_w];
assign v534ibus[data_w*4 +:data_w] = c920obus[data_w*0 +:data_w];
assign c920ibus[temp_w*1 +:temp_w] = v691obus[temp_w*4 +:temp_w];
assign v691ibus[data_w*4 +:data_w] = c920obus[data_w*1 +:data_w];
assign c920ibus[temp_w*2 +:temp_w] = v990obus[temp_w*2 +:temp_w];
assign v990ibus[data_w*2 +:data_w] = c920obus[data_w*2 +:data_w];
assign c920ibus[temp_w*3 +:temp_w] = v1088obus[temp_w*4 +:temp_w];
assign v1088ibus[data_w*4 +:data_w] = c920obus[data_w*3 +:data_w];
assign c920ibus[temp_w*4 +:temp_w] = v2072obus[temp_w*1 +:temp_w];
assign v2072ibus[data_w*1 +:data_w] = c920obus[data_w*4 +:data_w];
assign c920ibus[temp_w*5 +:temp_w] = v2168obus[temp_w*0 +:temp_w];
assign v2168ibus[data_w*0 +:data_w] = c920obus[data_w*5 +:data_w];
assign c921ibus[temp_w*0 +:temp_w] = v535obus[temp_w*4 +:temp_w];
assign v535ibus[data_w*4 +:data_w] = c921obus[data_w*0 +:data_w];
assign c921ibus[temp_w*1 +:temp_w] = v692obus[temp_w*4 +:temp_w];
assign v692ibus[data_w*4 +:data_w] = c921obus[data_w*1 +:data_w];
assign c921ibus[temp_w*2 +:temp_w] = v991obus[temp_w*2 +:temp_w];
assign v991ibus[data_w*2 +:data_w] = c921obus[data_w*2 +:data_w];
assign c921ibus[temp_w*3 +:temp_w] = v1089obus[temp_w*4 +:temp_w];
assign v1089ibus[data_w*4 +:data_w] = c921obus[data_w*3 +:data_w];
assign c921ibus[temp_w*4 +:temp_w] = v2073obus[temp_w*1 +:temp_w];
assign v2073ibus[data_w*1 +:data_w] = c921obus[data_w*4 +:data_w];
assign c921ibus[temp_w*5 +:temp_w] = v2169obus[temp_w*0 +:temp_w];
assign v2169ibus[data_w*0 +:data_w] = c921obus[data_w*5 +:data_w];
assign c922ibus[temp_w*0 +:temp_w] = v536obus[temp_w*4 +:temp_w];
assign v536ibus[data_w*4 +:data_w] = c922obus[data_w*0 +:data_w];
assign c922ibus[temp_w*1 +:temp_w] = v693obus[temp_w*4 +:temp_w];
assign v693ibus[data_w*4 +:data_w] = c922obus[data_w*1 +:data_w];
assign c922ibus[temp_w*2 +:temp_w] = v992obus[temp_w*2 +:temp_w];
assign v992ibus[data_w*2 +:data_w] = c922obus[data_w*2 +:data_w];
assign c922ibus[temp_w*3 +:temp_w] = v1090obus[temp_w*4 +:temp_w];
assign v1090ibus[data_w*4 +:data_w] = c922obus[data_w*3 +:data_w];
assign c922ibus[temp_w*4 +:temp_w] = v2074obus[temp_w*1 +:temp_w];
assign v2074ibus[data_w*1 +:data_w] = c922obus[data_w*4 +:data_w];
assign c922ibus[temp_w*5 +:temp_w] = v2170obus[temp_w*0 +:temp_w];
assign v2170ibus[data_w*0 +:data_w] = c922obus[data_w*5 +:data_w];
assign c923ibus[temp_w*0 +:temp_w] = v537obus[temp_w*4 +:temp_w];
assign v537ibus[data_w*4 +:data_w] = c923obus[data_w*0 +:data_w];
assign c923ibus[temp_w*1 +:temp_w] = v694obus[temp_w*4 +:temp_w];
assign v694ibus[data_w*4 +:data_w] = c923obus[data_w*1 +:data_w];
assign c923ibus[temp_w*2 +:temp_w] = v993obus[temp_w*2 +:temp_w];
assign v993ibus[data_w*2 +:data_w] = c923obus[data_w*2 +:data_w];
assign c923ibus[temp_w*3 +:temp_w] = v1091obus[temp_w*4 +:temp_w];
assign v1091ibus[data_w*4 +:data_w] = c923obus[data_w*3 +:data_w];
assign c923ibus[temp_w*4 +:temp_w] = v2075obus[temp_w*1 +:temp_w];
assign v2075ibus[data_w*1 +:data_w] = c923obus[data_w*4 +:data_w];
assign c923ibus[temp_w*5 +:temp_w] = v2171obus[temp_w*0 +:temp_w];
assign v2171ibus[data_w*0 +:data_w] = c923obus[data_w*5 +:data_w];
assign c924ibus[temp_w*0 +:temp_w] = v538obus[temp_w*4 +:temp_w];
assign v538ibus[data_w*4 +:data_w] = c924obus[data_w*0 +:data_w];
assign c924ibus[temp_w*1 +:temp_w] = v695obus[temp_w*4 +:temp_w];
assign v695ibus[data_w*4 +:data_w] = c924obus[data_w*1 +:data_w];
assign c924ibus[temp_w*2 +:temp_w] = v994obus[temp_w*2 +:temp_w];
assign v994ibus[data_w*2 +:data_w] = c924obus[data_w*2 +:data_w];
assign c924ibus[temp_w*3 +:temp_w] = v1092obus[temp_w*4 +:temp_w];
assign v1092ibus[data_w*4 +:data_w] = c924obus[data_w*3 +:data_w];
assign c924ibus[temp_w*4 +:temp_w] = v2076obus[temp_w*1 +:temp_w];
assign v2076ibus[data_w*1 +:data_w] = c924obus[data_w*4 +:data_w];
assign c924ibus[temp_w*5 +:temp_w] = v2172obus[temp_w*0 +:temp_w];
assign v2172ibus[data_w*0 +:data_w] = c924obus[data_w*5 +:data_w];
assign c925ibus[temp_w*0 +:temp_w] = v539obus[temp_w*4 +:temp_w];
assign v539ibus[data_w*4 +:data_w] = c925obus[data_w*0 +:data_w];
assign c925ibus[temp_w*1 +:temp_w] = v696obus[temp_w*4 +:temp_w];
assign v696ibus[data_w*4 +:data_w] = c925obus[data_w*1 +:data_w];
assign c925ibus[temp_w*2 +:temp_w] = v995obus[temp_w*2 +:temp_w];
assign v995ibus[data_w*2 +:data_w] = c925obus[data_w*2 +:data_w];
assign c925ibus[temp_w*3 +:temp_w] = v1093obus[temp_w*4 +:temp_w];
assign v1093ibus[data_w*4 +:data_w] = c925obus[data_w*3 +:data_w];
assign c925ibus[temp_w*4 +:temp_w] = v2077obus[temp_w*1 +:temp_w];
assign v2077ibus[data_w*1 +:data_w] = c925obus[data_w*4 +:data_w];
assign c925ibus[temp_w*5 +:temp_w] = v2173obus[temp_w*0 +:temp_w];
assign v2173ibus[data_w*0 +:data_w] = c925obus[data_w*5 +:data_w];
assign c926ibus[temp_w*0 +:temp_w] = v540obus[temp_w*4 +:temp_w];
assign v540ibus[data_w*4 +:data_w] = c926obus[data_w*0 +:data_w];
assign c926ibus[temp_w*1 +:temp_w] = v697obus[temp_w*4 +:temp_w];
assign v697ibus[data_w*4 +:data_w] = c926obus[data_w*1 +:data_w];
assign c926ibus[temp_w*2 +:temp_w] = v996obus[temp_w*2 +:temp_w];
assign v996ibus[data_w*2 +:data_w] = c926obus[data_w*2 +:data_w];
assign c926ibus[temp_w*3 +:temp_w] = v1094obus[temp_w*4 +:temp_w];
assign v1094ibus[data_w*4 +:data_w] = c926obus[data_w*3 +:data_w];
assign c926ibus[temp_w*4 +:temp_w] = v2078obus[temp_w*1 +:temp_w];
assign v2078ibus[data_w*1 +:data_w] = c926obus[data_w*4 +:data_w];
assign c926ibus[temp_w*5 +:temp_w] = v2174obus[temp_w*0 +:temp_w];
assign v2174ibus[data_w*0 +:data_w] = c926obus[data_w*5 +:data_w];
assign c927ibus[temp_w*0 +:temp_w] = v541obus[temp_w*4 +:temp_w];
assign v541ibus[data_w*4 +:data_w] = c927obus[data_w*0 +:data_w];
assign c927ibus[temp_w*1 +:temp_w] = v698obus[temp_w*4 +:temp_w];
assign v698ibus[data_w*4 +:data_w] = c927obus[data_w*1 +:data_w];
assign c927ibus[temp_w*2 +:temp_w] = v997obus[temp_w*2 +:temp_w];
assign v997ibus[data_w*2 +:data_w] = c927obus[data_w*2 +:data_w];
assign c927ibus[temp_w*3 +:temp_w] = v1095obus[temp_w*4 +:temp_w];
assign v1095ibus[data_w*4 +:data_w] = c927obus[data_w*3 +:data_w];
assign c927ibus[temp_w*4 +:temp_w] = v2079obus[temp_w*1 +:temp_w];
assign v2079ibus[data_w*1 +:data_w] = c927obus[data_w*4 +:data_w];
assign c927ibus[temp_w*5 +:temp_w] = v2175obus[temp_w*0 +:temp_w];
assign v2175ibus[data_w*0 +:data_w] = c927obus[data_w*5 +:data_w];
assign c928ibus[temp_w*0 +:temp_w] = v542obus[temp_w*4 +:temp_w];
assign v542ibus[data_w*4 +:data_w] = c928obus[data_w*0 +:data_w];
assign c928ibus[temp_w*1 +:temp_w] = v699obus[temp_w*4 +:temp_w];
assign v699ibus[data_w*4 +:data_w] = c928obus[data_w*1 +:data_w];
assign c928ibus[temp_w*2 +:temp_w] = v998obus[temp_w*2 +:temp_w];
assign v998ibus[data_w*2 +:data_w] = c928obus[data_w*2 +:data_w];
assign c928ibus[temp_w*3 +:temp_w] = v1096obus[temp_w*4 +:temp_w];
assign v1096ibus[data_w*4 +:data_w] = c928obus[data_w*3 +:data_w];
assign c928ibus[temp_w*4 +:temp_w] = v2080obus[temp_w*1 +:temp_w];
assign v2080ibus[data_w*1 +:data_w] = c928obus[data_w*4 +:data_w];
assign c928ibus[temp_w*5 +:temp_w] = v2176obus[temp_w*0 +:temp_w];
assign v2176ibus[data_w*0 +:data_w] = c928obus[data_w*5 +:data_w];
assign c929ibus[temp_w*0 +:temp_w] = v543obus[temp_w*4 +:temp_w];
assign v543ibus[data_w*4 +:data_w] = c929obus[data_w*0 +:data_w];
assign c929ibus[temp_w*1 +:temp_w] = v700obus[temp_w*4 +:temp_w];
assign v700ibus[data_w*4 +:data_w] = c929obus[data_w*1 +:data_w];
assign c929ibus[temp_w*2 +:temp_w] = v999obus[temp_w*2 +:temp_w];
assign v999ibus[data_w*2 +:data_w] = c929obus[data_w*2 +:data_w];
assign c929ibus[temp_w*3 +:temp_w] = v1097obus[temp_w*4 +:temp_w];
assign v1097ibus[data_w*4 +:data_w] = c929obus[data_w*3 +:data_w];
assign c929ibus[temp_w*4 +:temp_w] = v2081obus[temp_w*1 +:temp_w];
assign v2081ibus[data_w*1 +:data_w] = c929obus[data_w*4 +:data_w];
assign c929ibus[temp_w*5 +:temp_w] = v2177obus[temp_w*0 +:temp_w];
assign v2177ibus[data_w*0 +:data_w] = c929obus[data_w*5 +:data_w];
assign c930ibus[temp_w*0 +:temp_w] = v544obus[temp_w*4 +:temp_w];
assign v544ibus[data_w*4 +:data_w] = c930obus[data_w*0 +:data_w];
assign c930ibus[temp_w*1 +:temp_w] = v701obus[temp_w*4 +:temp_w];
assign v701ibus[data_w*4 +:data_w] = c930obus[data_w*1 +:data_w];
assign c930ibus[temp_w*2 +:temp_w] = v1000obus[temp_w*2 +:temp_w];
assign v1000ibus[data_w*2 +:data_w] = c930obus[data_w*2 +:data_w];
assign c930ibus[temp_w*3 +:temp_w] = v1098obus[temp_w*4 +:temp_w];
assign v1098ibus[data_w*4 +:data_w] = c930obus[data_w*3 +:data_w];
assign c930ibus[temp_w*4 +:temp_w] = v2082obus[temp_w*1 +:temp_w];
assign v2082ibus[data_w*1 +:data_w] = c930obus[data_w*4 +:data_w];
assign c930ibus[temp_w*5 +:temp_w] = v2178obus[temp_w*0 +:temp_w];
assign v2178ibus[data_w*0 +:data_w] = c930obus[data_w*5 +:data_w];
assign c931ibus[temp_w*0 +:temp_w] = v545obus[temp_w*4 +:temp_w];
assign v545ibus[data_w*4 +:data_w] = c931obus[data_w*0 +:data_w];
assign c931ibus[temp_w*1 +:temp_w] = v702obus[temp_w*4 +:temp_w];
assign v702ibus[data_w*4 +:data_w] = c931obus[data_w*1 +:data_w];
assign c931ibus[temp_w*2 +:temp_w] = v1001obus[temp_w*2 +:temp_w];
assign v1001ibus[data_w*2 +:data_w] = c931obus[data_w*2 +:data_w];
assign c931ibus[temp_w*3 +:temp_w] = v1099obus[temp_w*4 +:temp_w];
assign v1099ibus[data_w*4 +:data_w] = c931obus[data_w*3 +:data_w];
assign c931ibus[temp_w*4 +:temp_w] = v2083obus[temp_w*1 +:temp_w];
assign v2083ibus[data_w*1 +:data_w] = c931obus[data_w*4 +:data_w];
assign c931ibus[temp_w*5 +:temp_w] = v2179obus[temp_w*0 +:temp_w];
assign v2179ibus[data_w*0 +:data_w] = c931obus[data_w*5 +:data_w];
assign c932ibus[temp_w*0 +:temp_w] = v546obus[temp_w*4 +:temp_w];
assign v546ibus[data_w*4 +:data_w] = c932obus[data_w*0 +:data_w];
assign c932ibus[temp_w*1 +:temp_w] = v703obus[temp_w*4 +:temp_w];
assign v703ibus[data_w*4 +:data_w] = c932obus[data_w*1 +:data_w];
assign c932ibus[temp_w*2 +:temp_w] = v1002obus[temp_w*2 +:temp_w];
assign v1002ibus[data_w*2 +:data_w] = c932obus[data_w*2 +:data_w];
assign c932ibus[temp_w*3 +:temp_w] = v1100obus[temp_w*4 +:temp_w];
assign v1100ibus[data_w*4 +:data_w] = c932obus[data_w*3 +:data_w];
assign c932ibus[temp_w*4 +:temp_w] = v2084obus[temp_w*1 +:temp_w];
assign v2084ibus[data_w*1 +:data_w] = c932obus[data_w*4 +:data_w];
assign c932ibus[temp_w*5 +:temp_w] = v2180obus[temp_w*0 +:temp_w];
assign v2180ibus[data_w*0 +:data_w] = c932obus[data_w*5 +:data_w];
assign c933ibus[temp_w*0 +:temp_w] = v547obus[temp_w*4 +:temp_w];
assign v547ibus[data_w*4 +:data_w] = c933obus[data_w*0 +:data_w];
assign c933ibus[temp_w*1 +:temp_w] = v704obus[temp_w*4 +:temp_w];
assign v704ibus[data_w*4 +:data_w] = c933obus[data_w*1 +:data_w];
assign c933ibus[temp_w*2 +:temp_w] = v1003obus[temp_w*2 +:temp_w];
assign v1003ibus[data_w*2 +:data_w] = c933obus[data_w*2 +:data_w];
assign c933ibus[temp_w*3 +:temp_w] = v1101obus[temp_w*4 +:temp_w];
assign v1101ibus[data_w*4 +:data_w] = c933obus[data_w*3 +:data_w];
assign c933ibus[temp_w*4 +:temp_w] = v2085obus[temp_w*1 +:temp_w];
assign v2085ibus[data_w*1 +:data_w] = c933obus[data_w*4 +:data_w];
assign c933ibus[temp_w*5 +:temp_w] = v2181obus[temp_w*0 +:temp_w];
assign v2181ibus[data_w*0 +:data_w] = c933obus[data_w*5 +:data_w];
assign c934ibus[temp_w*0 +:temp_w] = v548obus[temp_w*4 +:temp_w];
assign v548ibus[data_w*4 +:data_w] = c934obus[data_w*0 +:data_w];
assign c934ibus[temp_w*1 +:temp_w] = v705obus[temp_w*4 +:temp_w];
assign v705ibus[data_w*4 +:data_w] = c934obus[data_w*1 +:data_w];
assign c934ibus[temp_w*2 +:temp_w] = v1004obus[temp_w*2 +:temp_w];
assign v1004ibus[data_w*2 +:data_w] = c934obus[data_w*2 +:data_w];
assign c934ibus[temp_w*3 +:temp_w] = v1102obus[temp_w*4 +:temp_w];
assign v1102ibus[data_w*4 +:data_w] = c934obus[data_w*3 +:data_w];
assign c934ibus[temp_w*4 +:temp_w] = v2086obus[temp_w*1 +:temp_w];
assign v2086ibus[data_w*1 +:data_w] = c934obus[data_w*4 +:data_w];
assign c934ibus[temp_w*5 +:temp_w] = v2182obus[temp_w*0 +:temp_w];
assign v2182ibus[data_w*0 +:data_w] = c934obus[data_w*5 +:data_w];
assign c935ibus[temp_w*0 +:temp_w] = v549obus[temp_w*4 +:temp_w];
assign v549ibus[data_w*4 +:data_w] = c935obus[data_w*0 +:data_w];
assign c935ibus[temp_w*1 +:temp_w] = v706obus[temp_w*4 +:temp_w];
assign v706ibus[data_w*4 +:data_w] = c935obus[data_w*1 +:data_w];
assign c935ibus[temp_w*2 +:temp_w] = v1005obus[temp_w*2 +:temp_w];
assign v1005ibus[data_w*2 +:data_w] = c935obus[data_w*2 +:data_w];
assign c935ibus[temp_w*3 +:temp_w] = v1103obus[temp_w*4 +:temp_w];
assign v1103ibus[data_w*4 +:data_w] = c935obus[data_w*3 +:data_w];
assign c935ibus[temp_w*4 +:temp_w] = v2087obus[temp_w*1 +:temp_w];
assign v2087ibus[data_w*1 +:data_w] = c935obus[data_w*4 +:data_w];
assign c935ibus[temp_w*5 +:temp_w] = v2183obus[temp_w*0 +:temp_w];
assign v2183ibus[data_w*0 +:data_w] = c935obus[data_w*5 +:data_w];
assign c936ibus[temp_w*0 +:temp_w] = v550obus[temp_w*4 +:temp_w];
assign v550ibus[data_w*4 +:data_w] = c936obus[data_w*0 +:data_w];
assign c936ibus[temp_w*1 +:temp_w] = v707obus[temp_w*4 +:temp_w];
assign v707ibus[data_w*4 +:data_w] = c936obus[data_w*1 +:data_w];
assign c936ibus[temp_w*2 +:temp_w] = v1006obus[temp_w*2 +:temp_w];
assign v1006ibus[data_w*2 +:data_w] = c936obus[data_w*2 +:data_w];
assign c936ibus[temp_w*3 +:temp_w] = v1104obus[temp_w*4 +:temp_w];
assign v1104ibus[data_w*4 +:data_w] = c936obus[data_w*3 +:data_w];
assign c936ibus[temp_w*4 +:temp_w] = v2088obus[temp_w*1 +:temp_w];
assign v2088ibus[data_w*1 +:data_w] = c936obus[data_w*4 +:data_w];
assign c936ibus[temp_w*5 +:temp_w] = v2184obus[temp_w*0 +:temp_w];
assign v2184ibus[data_w*0 +:data_w] = c936obus[data_w*5 +:data_w];
assign c937ibus[temp_w*0 +:temp_w] = v551obus[temp_w*4 +:temp_w];
assign v551ibus[data_w*4 +:data_w] = c937obus[data_w*0 +:data_w];
assign c937ibus[temp_w*1 +:temp_w] = v708obus[temp_w*4 +:temp_w];
assign v708ibus[data_w*4 +:data_w] = c937obus[data_w*1 +:data_w];
assign c937ibus[temp_w*2 +:temp_w] = v1007obus[temp_w*2 +:temp_w];
assign v1007ibus[data_w*2 +:data_w] = c937obus[data_w*2 +:data_w];
assign c937ibus[temp_w*3 +:temp_w] = v1105obus[temp_w*4 +:temp_w];
assign v1105ibus[data_w*4 +:data_w] = c937obus[data_w*3 +:data_w];
assign c937ibus[temp_w*4 +:temp_w] = v2089obus[temp_w*1 +:temp_w];
assign v2089ibus[data_w*1 +:data_w] = c937obus[data_w*4 +:data_w];
assign c937ibus[temp_w*5 +:temp_w] = v2185obus[temp_w*0 +:temp_w];
assign v2185ibus[data_w*0 +:data_w] = c937obus[data_w*5 +:data_w];
assign c938ibus[temp_w*0 +:temp_w] = v552obus[temp_w*4 +:temp_w];
assign v552ibus[data_w*4 +:data_w] = c938obus[data_w*0 +:data_w];
assign c938ibus[temp_w*1 +:temp_w] = v709obus[temp_w*4 +:temp_w];
assign v709ibus[data_w*4 +:data_w] = c938obus[data_w*1 +:data_w];
assign c938ibus[temp_w*2 +:temp_w] = v1008obus[temp_w*2 +:temp_w];
assign v1008ibus[data_w*2 +:data_w] = c938obus[data_w*2 +:data_w];
assign c938ibus[temp_w*3 +:temp_w] = v1106obus[temp_w*4 +:temp_w];
assign v1106ibus[data_w*4 +:data_w] = c938obus[data_w*3 +:data_w];
assign c938ibus[temp_w*4 +:temp_w] = v2090obus[temp_w*1 +:temp_w];
assign v2090ibus[data_w*1 +:data_w] = c938obus[data_w*4 +:data_w];
assign c938ibus[temp_w*5 +:temp_w] = v2186obus[temp_w*0 +:temp_w];
assign v2186ibus[data_w*0 +:data_w] = c938obus[data_w*5 +:data_w];
assign c939ibus[temp_w*0 +:temp_w] = v553obus[temp_w*4 +:temp_w];
assign v553ibus[data_w*4 +:data_w] = c939obus[data_w*0 +:data_w];
assign c939ibus[temp_w*1 +:temp_w] = v710obus[temp_w*4 +:temp_w];
assign v710ibus[data_w*4 +:data_w] = c939obus[data_w*1 +:data_w];
assign c939ibus[temp_w*2 +:temp_w] = v1009obus[temp_w*2 +:temp_w];
assign v1009ibus[data_w*2 +:data_w] = c939obus[data_w*2 +:data_w];
assign c939ibus[temp_w*3 +:temp_w] = v1107obus[temp_w*4 +:temp_w];
assign v1107ibus[data_w*4 +:data_w] = c939obus[data_w*3 +:data_w];
assign c939ibus[temp_w*4 +:temp_w] = v2091obus[temp_w*1 +:temp_w];
assign v2091ibus[data_w*1 +:data_w] = c939obus[data_w*4 +:data_w];
assign c939ibus[temp_w*5 +:temp_w] = v2187obus[temp_w*0 +:temp_w];
assign v2187ibus[data_w*0 +:data_w] = c939obus[data_w*5 +:data_w];
assign c940ibus[temp_w*0 +:temp_w] = v554obus[temp_w*4 +:temp_w];
assign v554ibus[data_w*4 +:data_w] = c940obus[data_w*0 +:data_w];
assign c940ibus[temp_w*1 +:temp_w] = v711obus[temp_w*4 +:temp_w];
assign v711ibus[data_w*4 +:data_w] = c940obus[data_w*1 +:data_w];
assign c940ibus[temp_w*2 +:temp_w] = v1010obus[temp_w*2 +:temp_w];
assign v1010ibus[data_w*2 +:data_w] = c940obus[data_w*2 +:data_w];
assign c940ibus[temp_w*3 +:temp_w] = v1108obus[temp_w*4 +:temp_w];
assign v1108ibus[data_w*4 +:data_w] = c940obus[data_w*3 +:data_w];
assign c940ibus[temp_w*4 +:temp_w] = v2092obus[temp_w*1 +:temp_w];
assign v2092ibus[data_w*1 +:data_w] = c940obus[data_w*4 +:data_w];
assign c940ibus[temp_w*5 +:temp_w] = v2188obus[temp_w*0 +:temp_w];
assign v2188ibus[data_w*0 +:data_w] = c940obus[data_w*5 +:data_w];
assign c941ibus[temp_w*0 +:temp_w] = v555obus[temp_w*4 +:temp_w];
assign v555ibus[data_w*4 +:data_w] = c941obus[data_w*0 +:data_w];
assign c941ibus[temp_w*1 +:temp_w] = v712obus[temp_w*4 +:temp_w];
assign v712ibus[data_w*4 +:data_w] = c941obus[data_w*1 +:data_w];
assign c941ibus[temp_w*2 +:temp_w] = v1011obus[temp_w*2 +:temp_w];
assign v1011ibus[data_w*2 +:data_w] = c941obus[data_w*2 +:data_w];
assign c941ibus[temp_w*3 +:temp_w] = v1109obus[temp_w*4 +:temp_w];
assign v1109ibus[data_w*4 +:data_w] = c941obus[data_w*3 +:data_w];
assign c941ibus[temp_w*4 +:temp_w] = v2093obus[temp_w*1 +:temp_w];
assign v2093ibus[data_w*1 +:data_w] = c941obus[data_w*4 +:data_w];
assign c941ibus[temp_w*5 +:temp_w] = v2189obus[temp_w*0 +:temp_w];
assign v2189ibus[data_w*0 +:data_w] = c941obus[data_w*5 +:data_w];
assign c942ibus[temp_w*0 +:temp_w] = v556obus[temp_w*4 +:temp_w];
assign v556ibus[data_w*4 +:data_w] = c942obus[data_w*0 +:data_w];
assign c942ibus[temp_w*1 +:temp_w] = v713obus[temp_w*4 +:temp_w];
assign v713ibus[data_w*4 +:data_w] = c942obus[data_w*1 +:data_w];
assign c942ibus[temp_w*2 +:temp_w] = v1012obus[temp_w*2 +:temp_w];
assign v1012ibus[data_w*2 +:data_w] = c942obus[data_w*2 +:data_w];
assign c942ibus[temp_w*3 +:temp_w] = v1110obus[temp_w*4 +:temp_w];
assign v1110ibus[data_w*4 +:data_w] = c942obus[data_w*3 +:data_w];
assign c942ibus[temp_w*4 +:temp_w] = v2094obus[temp_w*1 +:temp_w];
assign v2094ibus[data_w*1 +:data_w] = c942obus[data_w*4 +:data_w];
assign c942ibus[temp_w*5 +:temp_w] = v2190obus[temp_w*0 +:temp_w];
assign v2190ibus[data_w*0 +:data_w] = c942obus[data_w*5 +:data_w];
assign c943ibus[temp_w*0 +:temp_w] = v557obus[temp_w*4 +:temp_w];
assign v557ibus[data_w*4 +:data_w] = c943obus[data_w*0 +:data_w];
assign c943ibus[temp_w*1 +:temp_w] = v714obus[temp_w*4 +:temp_w];
assign v714ibus[data_w*4 +:data_w] = c943obus[data_w*1 +:data_w];
assign c943ibus[temp_w*2 +:temp_w] = v1013obus[temp_w*2 +:temp_w];
assign v1013ibus[data_w*2 +:data_w] = c943obus[data_w*2 +:data_w];
assign c943ibus[temp_w*3 +:temp_w] = v1111obus[temp_w*4 +:temp_w];
assign v1111ibus[data_w*4 +:data_w] = c943obus[data_w*3 +:data_w];
assign c943ibus[temp_w*4 +:temp_w] = v2095obus[temp_w*1 +:temp_w];
assign v2095ibus[data_w*1 +:data_w] = c943obus[data_w*4 +:data_w];
assign c943ibus[temp_w*5 +:temp_w] = v2191obus[temp_w*0 +:temp_w];
assign v2191ibus[data_w*0 +:data_w] = c943obus[data_w*5 +:data_w];
assign c944ibus[temp_w*0 +:temp_w] = v558obus[temp_w*4 +:temp_w];
assign v558ibus[data_w*4 +:data_w] = c944obus[data_w*0 +:data_w];
assign c944ibus[temp_w*1 +:temp_w] = v715obus[temp_w*4 +:temp_w];
assign v715ibus[data_w*4 +:data_w] = c944obus[data_w*1 +:data_w];
assign c944ibus[temp_w*2 +:temp_w] = v1014obus[temp_w*2 +:temp_w];
assign v1014ibus[data_w*2 +:data_w] = c944obus[data_w*2 +:data_w];
assign c944ibus[temp_w*3 +:temp_w] = v1112obus[temp_w*4 +:temp_w];
assign v1112ibus[data_w*4 +:data_w] = c944obus[data_w*3 +:data_w];
assign c944ibus[temp_w*4 +:temp_w] = v2096obus[temp_w*1 +:temp_w];
assign v2096ibus[data_w*1 +:data_w] = c944obus[data_w*4 +:data_w];
assign c944ibus[temp_w*5 +:temp_w] = v2192obus[temp_w*0 +:temp_w];
assign v2192ibus[data_w*0 +:data_w] = c944obus[data_w*5 +:data_w];
assign c945ibus[temp_w*0 +:temp_w] = v559obus[temp_w*4 +:temp_w];
assign v559ibus[data_w*4 +:data_w] = c945obus[data_w*0 +:data_w];
assign c945ibus[temp_w*1 +:temp_w] = v716obus[temp_w*4 +:temp_w];
assign v716ibus[data_w*4 +:data_w] = c945obus[data_w*1 +:data_w];
assign c945ibus[temp_w*2 +:temp_w] = v1015obus[temp_w*2 +:temp_w];
assign v1015ibus[data_w*2 +:data_w] = c945obus[data_w*2 +:data_w];
assign c945ibus[temp_w*3 +:temp_w] = v1113obus[temp_w*4 +:temp_w];
assign v1113ibus[data_w*4 +:data_w] = c945obus[data_w*3 +:data_w];
assign c945ibus[temp_w*4 +:temp_w] = v2097obus[temp_w*1 +:temp_w];
assign v2097ibus[data_w*1 +:data_w] = c945obus[data_w*4 +:data_w];
assign c945ibus[temp_w*5 +:temp_w] = v2193obus[temp_w*0 +:temp_w];
assign v2193ibus[data_w*0 +:data_w] = c945obus[data_w*5 +:data_w];
assign c946ibus[temp_w*0 +:temp_w] = v560obus[temp_w*4 +:temp_w];
assign v560ibus[data_w*4 +:data_w] = c946obus[data_w*0 +:data_w];
assign c946ibus[temp_w*1 +:temp_w] = v717obus[temp_w*4 +:temp_w];
assign v717ibus[data_w*4 +:data_w] = c946obus[data_w*1 +:data_w];
assign c946ibus[temp_w*2 +:temp_w] = v1016obus[temp_w*2 +:temp_w];
assign v1016ibus[data_w*2 +:data_w] = c946obus[data_w*2 +:data_w];
assign c946ibus[temp_w*3 +:temp_w] = v1114obus[temp_w*4 +:temp_w];
assign v1114ibus[data_w*4 +:data_w] = c946obus[data_w*3 +:data_w];
assign c946ibus[temp_w*4 +:temp_w] = v2098obus[temp_w*1 +:temp_w];
assign v2098ibus[data_w*1 +:data_w] = c946obus[data_w*4 +:data_w];
assign c946ibus[temp_w*5 +:temp_w] = v2194obus[temp_w*0 +:temp_w];
assign v2194ibus[data_w*0 +:data_w] = c946obus[data_w*5 +:data_w];
assign c947ibus[temp_w*0 +:temp_w] = v561obus[temp_w*4 +:temp_w];
assign v561ibus[data_w*4 +:data_w] = c947obus[data_w*0 +:data_w];
assign c947ibus[temp_w*1 +:temp_w] = v718obus[temp_w*4 +:temp_w];
assign v718ibus[data_w*4 +:data_w] = c947obus[data_w*1 +:data_w];
assign c947ibus[temp_w*2 +:temp_w] = v1017obus[temp_w*2 +:temp_w];
assign v1017ibus[data_w*2 +:data_w] = c947obus[data_w*2 +:data_w];
assign c947ibus[temp_w*3 +:temp_w] = v1115obus[temp_w*4 +:temp_w];
assign v1115ibus[data_w*4 +:data_w] = c947obus[data_w*3 +:data_w];
assign c947ibus[temp_w*4 +:temp_w] = v2099obus[temp_w*1 +:temp_w];
assign v2099ibus[data_w*1 +:data_w] = c947obus[data_w*4 +:data_w];
assign c947ibus[temp_w*5 +:temp_w] = v2195obus[temp_w*0 +:temp_w];
assign v2195ibus[data_w*0 +:data_w] = c947obus[data_w*5 +:data_w];
assign c948ibus[temp_w*0 +:temp_w] = v562obus[temp_w*4 +:temp_w];
assign v562ibus[data_w*4 +:data_w] = c948obus[data_w*0 +:data_w];
assign c948ibus[temp_w*1 +:temp_w] = v719obus[temp_w*4 +:temp_w];
assign v719ibus[data_w*4 +:data_w] = c948obus[data_w*1 +:data_w];
assign c948ibus[temp_w*2 +:temp_w] = v1018obus[temp_w*2 +:temp_w];
assign v1018ibus[data_w*2 +:data_w] = c948obus[data_w*2 +:data_w];
assign c948ibus[temp_w*3 +:temp_w] = v1116obus[temp_w*4 +:temp_w];
assign v1116ibus[data_w*4 +:data_w] = c948obus[data_w*3 +:data_w];
assign c948ibus[temp_w*4 +:temp_w] = v2100obus[temp_w*1 +:temp_w];
assign v2100ibus[data_w*1 +:data_w] = c948obus[data_w*4 +:data_w];
assign c948ibus[temp_w*5 +:temp_w] = v2196obus[temp_w*0 +:temp_w];
assign v2196ibus[data_w*0 +:data_w] = c948obus[data_w*5 +:data_w];
assign c949ibus[temp_w*0 +:temp_w] = v563obus[temp_w*4 +:temp_w];
assign v563ibus[data_w*4 +:data_w] = c949obus[data_w*0 +:data_w];
assign c949ibus[temp_w*1 +:temp_w] = v720obus[temp_w*4 +:temp_w];
assign v720ibus[data_w*4 +:data_w] = c949obus[data_w*1 +:data_w];
assign c949ibus[temp_w*2 +:temp_w] = v1019obus[temp_w*2 +:temp_w];
assign v1019ibus[data_w*2 +:data_w] = c949obus[data_w*2 +:data_w];
assign c949ibus[temp_w*3 +:temp_w] = v1117obus[temp_w*4 +:temp_w];
assign v1117ibus[data_w*4 +:data_w] = c949obus[data_w*3 +:data_w];
assign c949ibus[temp_w*4 +:temp_w] = v2101obus[temp_w*1 +:temp_w];
assign v2101ibus[data_w*1 +:data_w] = c949obus[data_w*4 +:data_w];
assign c949ibus[temp_w*5 +:temp_w] = v2197obus[temp_w*0 +:temp_w];
assign v2197ibus[data_w*0 +:data_w] = c949obus[data_w*5 +:data_w];
assign c950ibus[temp_w*0 +:temp_w] = v564obus[temp_w*4 +:temp_w];
assign v564ibus[data_w*4 +:data_w] = c950obus[data_w*0 +:data_w];
assign c950ibus[temp_w*1 +:temp_w] = v721obus[temp_w*4 +:temp_w];
assign v721ibus[data_w*4 +:data_w] = c950obus[data_w*1 +:data_w];
assign c950ibus[temp_w*2 +:temp_w] = v1020obus[temp_w*2 +:temp_w];
assign v1020ibus[data_w*2 +:data_w] = c950obus[data_w*2 +:data_w];
assign c950ibus[temp_w*3 +:temp_w] = v1118obus[temp_w*4 +:temp_w];
assign v1118ibus[data_w*4 +:data_w] = c950obus[data_w*3 +:data_w];
assign c950ibus[temp_w*4 +:temp_w] = v2102obus[temp_w*1 +:temp_w];
assign v2102ibus[data_w*1 +:data_w] = c950obus[data_w*4 +:data_w];
assign c950ibus[temp_w*5 +:temp_w] = v2198obus[temp_w*0 +:temp_w];
assign v2198ibus[data_w*0 +:data_w] = c950obus[data_w*5 +:data_w];
assign c951ibus[temp_w*0 +:temp_w] = v565obus[temp_w*4 +:temp_w];
assign v565ibus[data_w*4 +:data_w] = c951obus[data_w*0 +:data_w];
assign c951ibus[temp_w*1 +:temp_w] = v722obus[temp_w*4 +:temp_w];
assign v722ibus[data_w*4 +:data_w] = c951obus[data_w*1 +:data_w];
assign c951ibus[temp_w*2 +:temp_w] = v1021obus[temp_w*2 +:temp_w];
assign v1021ibus[data_w*2 +:data_w] = c951obus[data_w*2 +:data_w];
assign c951ibus[temp_w*3 +:temp_w] = v1119obus[temp_w*4 +:temp_w];
assign v1119ibus[data_w*4 +:data_w] = c951obus[data_w*3 +:data_w];
assign c951ibus[temp_w*4 +:temp_w] = v2103obus[temp_w*1 +:temp_w];
assign v2103ibus[data_w*1 +:data_w] = c951obus[data_w*4 +:data_w];
assign c951ibus[temp_w*5 +:temp_w] = v2199obus[temp_w*0 +:temp_w];
assign v2199ibus[data_w*0 +:data_w] = c951obus[data_w*5 +:data_w];
assign c952ibus[temp_w*0 +:temp_w] = v566obus[temp_w*4 +:temp_w];
assign v566ibus[data_w*4 +:data_w] = c952obus[data_w*0 +:data_w];
assign c952ibus[temp_w*1 +:temp_w] = v723obus[temp_w*4 +:temp_w];
assign v723ibus[data_w*4 +:data_w] = c952obus[data_w*1 +:data_w];
assign c952ibus[temp_w*2 +:temp_w] = v1022obus[temp_w*2 +:temp_w];
assign v1022ibus[data_w*2 +:data_w] = c952obus[data_w*2 +:data_w];
assign c952ibus[temp_w*3 +:temp_w] = v1120obus[temp_w*4 +:temp_w];
assign v1120ibus[data_w*4 +:data_w] = c952obus[data_w*3 +:data_w];
assign c952ibus[temp_w*4 +:temp_w] = v2104obus[temp_w*1 +:temp_w];
assign v2104ibus[data_w*1 +:data_w] = c952obus[data_w*4 +:data_w];
assign c952ibus[temp_w*5 +:temp_w] = v2200obus[temp_w*0 +:temp_w];
assign v2200ibus[data_w*0 +:data_w] = c952obus[data_w*5 +:data_w];
assign c953ibus[temp_w*0 +:temp_w] = v567obus[temp_w*4 +:temp_w];
assign v567ibus[data_w*4 +:data_w] = c953obus[data_w*0 +:data_w];
assign c953ibus[temp_w*1 +:temp_w] = v724obus[temp_w*4 +:temp_w];
assign v724ibus[data_w*4 +:data_w] = c953obus[data_w*1 +:data_w];
assign c953ibus[temp_w*2 +:temp_w] = v1023obus[temp_w*2 +:temp_w];
assign v1023ibus[data_w*2 +:data_w] = c953obus[data_w*2 +:data_w];
assign c953ibus[temp_w*3 +:temp_w] = v1121obus[temp_w*4 +:temp_w];
assign v1121ibus[data_w*4 +:data_w] = c953obus[data_w*3 +:data_w];
assign c953ibus[temp_w*4 +:temp_w] = v2105obus[temp_w*1 +:temp_w];
assign v2105ibus[data_w*1 +:data_w] = c953obus[data_w*4 +:data_w];
assign c953ibus[temp_w*5 +:temp_w] = v2201obus[temp_w*0 +:temp_w];
assign v2201ibus[data_w*0 +:data_w] = c953obus[data_w*5 +:data_w];
assign c954ibus[temp_w*0 +:temp_w] = v568obus[temp_w*4 +:temp_w];
assign v568ibus[data_w*4 +:data_w] = c954obus[data_w*0 +:data_w];
assign c954ibus[temp_w*1 +:temp_w] = v725obus[temp_w*4 +:temp_w];
assign v725ibus[data_w*4 +:data_w] = c954obus[data_w*1 +:data_w];
assign c954ibus[temp_w*2 +:temp_w] = v1024obus[temp_w*2 +:temp_w];
assign v1024ibus[data_w*2 +:data_w] = c954obus[data_w*2 +:data_w];
assign c954ibus[temp_w*3 +:temp_w] = v1122obus[temp_w*4 +:temp_w];
assign v1122ibus[data_w*4 +:data_w] = c954obus[data_w*3 +:data_w];
assign c954ibus[temp_w*4 +:temp_w] = v2106obus[temp_w*1 +:temp_w];
assign v2106ibus[data_w*1 +:data_w] = c954obus[data_w*4 +:data_w];
assign c954ibus[temp_w*5 +:temp_w] = v2202obus[temp_w*0 +:temp_w];
assign v2202ibus[data_w*0 +:data_w] = c954obus[data_w*5 +:data_w];
assign c955ibus[temp_w*0 +:temp_w] = v569obus[temp_w*4 +:temp_w];
assign v569ibus[data_w*4 +:data_w] = c955obus[data_w*0 +:data_w];
assign c955ibus[temp_w*1 +:temp_w] = v726obus[temp_w*4 +:temp_w];
assign v726ibus[data_w*4 +:data_w] = c955obus[data_w*1 +:data_w];
assign c955ibus[temp_w*2 +:temp_w] = v1025obus[temp_w*2 +:temp_w];
assign v1025ibus[data_w*2 +:data_w] = c955obus[data_w*2 +:data_w];
assign c955ibus[temp_w*3 +:temp_w] = v1123obus[temp_w*4 +:temp_w];
assign v1123ibus[data_w*4 +:data_w] = c955obus[data_w*3 +:data_w];
assign c955ibus[temp_w*4 +:temp_w] = v2107obus[temp_w*1 +:temp_w];
assign v2107ibus[data_w*1 +:data_w] = c955obus[data_w*4 +:data_w];
assign c955ibus[temp_w*5 +:temp_w] = v2203obus[temp_w*0 +:temp_w];
assign v2203ibus[data_w*0 +:data_w] = c955obus[data_w*5 +:data_w];
assign c956ibus[temp_w*0 +:temp_w] = v570obus[temp_w*4 +:temp_w];
assign v570ibus[data_w*4 +:data_w] = c956obus[data_w*0 +:data_w];
assign c956ibus[temp_w*1 +:temp_w] = v727obus[temp_w*4 +:temp_w];
assign v727ibus[data_w*4 +:data_w] = c956obus[data_w*1 +:data_w];
assign c956ibus[temp_w*2 +:temp_w] = v1026obus[temp_w*2 +:temp_w];
assign v1026ibus[data_w*2 +:data_w] = c956obus[data_w*2 +:data_w];
assign c956ibus[temp_w*3 +:temp_w] = v1124obus[temp_w*4 +:temp_w];
assign v1124ibus[data_w*4 +:data_w] = c956obus[data_w*3 +:data_w];
assign c956ibus[temp_w*4 +:temp_w] = v2108obus[temp_w*1 +:temp_w];
assign v2108ibus[data_w*1 +:data_w] = c956obus[data_w*4 +:data_w];
assign c956ibus[temp_w*5 +:temp_w] = v2204obus[temp_w*0 +:temp_w];
assign v2204ibus[data_w*0 +:data_w] = c956obus[data_w*5 +:data_w];
assign c957ibus[temp_w*0 +:temp_w] = v571obus[temp_w*4 +:temp_w];
assign v571ibus[data_w*4 +:data_w] = c957obus[data_w*0 +:data_w];
assign c957ibus[temp_w*1 +:temp_w] = v728obus[temp_w*4 +:temp_w];
assign v728ibus[data_w*4 +:data_w] = c957obus[data_w*1 +:data_w];
assign c957ibus[temp_w*2 +:temp_w] = v1027obus[temp_w*2 +:temp_w];
assign v1027ibus[data_w*2 +:data_w] = c957obus[data_w*2 +:data_w];
assign c957ibus[temp_w*3 +:temp_w] = v1125obus[temp_w*4 +:temp_w];
assign v1125ibus[data_w*4 +:data_w] = c957obus[data_w*3 +:data_w];
assign c957ibus[temp_w*4 +:temp_w] = v2109obus[temp_w*1 +:temp_w];
assign v2109ibus[data_w*1 +:data_w] = c957obus[data_w*4 +:data_w];
assign c957ibus[temp_w*5 +:temp_w] = v2205obus[temp_w*0 +:temp_w];
assign v2205ibus[data_w*0 +:data_w] = c957obus[data_w*5 +:data_w];
assign c958ibus[temp_w*0 +:temp_w] = v572obus[temp_w*4 +:temp_w];
assign v572ibus[data_w*4 +:data_w] = c958obus[data_w*0 +:data_w];
assign c958ibus[temp_w*1 +:temp_w] = v729obus[temp_w*4 +:temp_w];
assign v729ibus[data_w*4 +:data_w] = c958obus[data_w*1 +:data_w];
assign c958ibus[temp_w*2 +:temp_w] = v1028obus[temp_w*2 +:temp_w];
assign v1028ibus[data_w*2 +:data_w] = c958obus[data_w*2 +:data_w];
assign c958ibus[temp_w*3 +:temp_w] = v1126obus[temp_w*4 +:temp_w];
assign v1126ibus[data_w*4 +:data_w] = c958obus[data_w*3 +:data_w];
assign c958ibus[temp_w*4 +:temp_w] = v2110obus[temp_w*1 +:temp_w];
assign v2110ibus[data_w*1 +:data_w] = c958obus[data_w*4 +:data_w];
assign c958ibus[temp_w*5 +:temp_w] = v2206obus[temp_w*0 +:temp_w];
assign v2206ibus[data_w*0 +:data_w] = c958obus[data_w*5 +:data_w];
assign c959ibus[temp_w*0 +:temp_w] = v573obus[temp_w*4 +:temp_w];
assign v573ibus[data_w*4 +:data_w] = c959obus[data_w*0 +:data_w];
assign c959ibus[temp_w*1 +:temp_w] = v730obus[temp_w*4 +:temp_w];
assign v730ibus[data_w*4 +:data_w] = c959obus[data_w*1 +:data_w];
assign c959ibus[temp_w*2 +:temp_w] = v1029obus[temp_w*2 +:temp_w];
assign v1029ibus[data_w*2 +:data_w] = c959obus[data_w*2 +:data_w];
assign c959ibus[temp_w*3 +:temp_w] = v1127obus[temp_w*4 +:temp_w];
assign v1127ibus[data_w*4 +:data_w] = c959obus[data_w*3 +:data_w];
assign c959ibus[temp_w*4 +:temp_w] = v2111obus[temp_w*1 +:temp_w];
assign v2111ibus[data_w*1 +:data_w] = c959obus[data_w*4 +:data_w];
assign c959ibus[temp_w*5 +:temp_w] = v2207obus[temp_w*0 +:temp_w];
assign v2207ibus[data_w*0 +:data_w] = c959obus[data_w*5 +:data_w];
assign c960ibus[temp_w*0 +:temp_w] = v199obus[temp_w*5 +:temp_w];
assign v199ibus[data_w*5 +:data_w] = c960obus[data_w*0 +:data_w];
assign c960ibus[temp_w*1 +:temp_w] = v353obus[temp_w*2 +:temp_w];
assign v353ibus[data_w*2 +:data_w] = c960obus[data_w*1 +:data_w];
assign c960ibus[temp_w*2 +:temp_w] = v807obus[temp_w*2 +:temp_w];
assign v807ibus[data_w*2 +:data_w] = c960obus[data_w*2 +:data_w];
assign c960ibus[temp_w*3 +:temp_w] = v913obus[temp_w*5 +:temp_w];
assign v913ibus[data_w*5 +:data_w] = c960obus[data_w*3 +:data_w];
assign c960ibus[temp_w*4 +:temp_w] = v2112obus[temp_w*1 +:temp_w];
assign v2112ibus[data_w*1 +:data_w] = c960obus[data_w*4 +:data_w];
assign c960ibus[temp_w*5 +:temp_w] = v2208obus[temp_w*0 +:temp_w];
assign v2208ibus[data_w*0 +:data_w] = c960obus[data_w*5 +:data_w];
assign c961ibus[temp_w*0 +:temp_w] = v200obus[temp_w*5 +:temp_w];
assign v200ibus[data_w*5 +:data_w] = c961obus[data_w*0 +:data_w];
assign c961ibus[temp_w*1 +:temp_w] = v354obus[temp_w*2 +:temp_w];
assign v354ibus[data_w*2 +:data_w] = c961obus[data_w*1 +:data_w];
assign c961ibus[temp_w*2 +:temp_w] = v808obus[temp_w*2 +:temp_w];
assign v808ibus[data_w*2 +:data_w] = c961obus[data_w*2 +:data_w];
assign c961ibus[temp_w*3 +:temp_w] = v914obus[temp_w*5 +:temp_w];
assign v914ibus[data_w*5 +:data_w] = c961obus[data_w*3 +:data_w];
assign c961ibus[temp_w*4 +:temp_w] = v2113obus[temp_w*1 +:temp_w];
assign v2113ibus[data_w*1 +:data_w] = c961obus[data_w*4 +:data_w];
assign c961ibus[temp_w*5 +:temp_w] = v2209obus[temp_w*0 +:temp_w];
assign v2209ibus[data_w*0 +:data_w] = c961obus[data_w*5 +:data_w];
assign c962ibus[temp_w*0 +:temp_w] = v201obus[temp_w*5 +:temp_w];
assign v201ibus[data_w*5 +:data_w] = c962obus[data_w*0 +:data_w];
assign c962ibus[temp_w*1 +:temp_w] = v355obus[temp_w*2 +:temp_w];
assign v355ibus[data_w*2 +:data_w] = c962obus[data_w*1 +:data_w];
assign c962ibus[temp_w*2 +:temp_w] = v809obus[temp_w*2 +:temp_w];
assign v809ibus[data_w*2 +:data_w] = c962obus[data_w*2 +:data_w];
assign c962ibus[temp_w*3 +:temp_w] = v915obus[temp_w*5 +:temp_w];
assign v915ibus[data_w*5 +:data_w] = c962obus[data_w*3 +:data_w];
assign c962ibus[temp_w*4 +:temp_w] = v2114obus[temp_w*1 +:temp_w];
assign v2114ibus[data_w*1 +:data_w] = c962obus[data_w*4 +:data_w];
assign c962ibus[temp_w*5 +:temp_w] = v2210obus[temp_w*0 +:temp_w];
assign v2210ibus[data_w*0 +:data_w] = c962obus[data_w*5 +:data_w];
assign c963ibus[temp_w*0 +:temp_w] = v202obus[temp_w*5 +:temp_w];
assign v202ibus[data_w*5 +:data_w] = c963obus[data_w*0 +:data_w];
assign c963ibus[temp_w*1 +:temp_w] = v356obus[temp_w*2 +:temp_w];
assign v356ibus[data_w*2 +:data_w] = c963obus[data_w*1 +:data_w];
assign c963ibus[temp_w*2 +:temp_w] = v810obus[temp_w*2 +:temp_w];
assign v810ibus[data_w*2 +:data_w] = c963obus[data_w*2 +:data_w];
assign c963ibus[temp_w*3 +:temp_w] = v916obus[temp_w*5 +:temp_w];
assign v916ibus[data_w*5 +:data_w] = c963obus[data_w*3 +:data_w];
assign c963ibus[temp_w*4 +:temp_w] = v2115obus[temp_w*1 +:temp_w];
assign v2115ibus[data_w*1 +:data_w] = c963obus[data_w*4 +:data_w];
assign c963ibus[temp_w*5 +:temp_w] = v2211obus[temp_w*0 +:temp_w];
assign v2211ibus[data_w*0 +:data_w] = c963obus[data_w*5 +:data_w];
assign c964ibus[temp_w*0 +:temp_w] = v203obus[temp_w*5 +:temp_w];
assign v203ibus[data_w*5 +:data_w] = c964obus[data_w*0 +:data_w];
assign c964ibus[temp_w*1 +:temp_w] = v357obus[temp_w*2 +:temp_w];
assign v357ibus[data_w*2 +:data_w] = c964obus[data_w*1 +:data_w];
assign c964ibus[temp_w*2 +:temp_w] = v811obus[temp_w*2 +:temp_w];
assign v811ibus[data_w*2 +:data_w] = c964obus[data_w*2 +:data_w];
assign c964ibus[temp_w*3 +:temp_w] = v917obus[temp_w*5 +:temp_w];
assign v917ibus[data_w*5 +:data_w] = c964obus[data_w*3 +:data_w];
assign c964ibus[temp_w*4 +:temp_w] = v2116obus[temp_w*1 +:temp_w];
assign v2116ibus[data_w*1 +:data_w] = c964obus[data_w*4 +:data_w];
assign c964ibus[temp_w*5 +:temp_w] = v2212obus[temp_w*0 +:temp_w];
assign v2212ibus[data_w*0 +:data_w] = c964obus[data_w*5 +:data_w];
assign c965ibus[temp_w*0 +:temp_w] = v204obus[temp_w*5 +:temp_w];
assign v204ibus[data_w*5 +:data_w] = c965obus[data_w*0 +:data_w];
assign c965ibus[temp_w*1 +:temp_w] = v358obus[temp_w*2 +:temp_w];
assign v358ibus[data_w*2 +:data_w] = c965obus[data_w*1 +:data_w];
assign c965ibus[temp_w*2 +:temp_w] = v812obus[temp_w*2 +:temp_w];
assign v812ibus[data_w*2 +:data_w] = c965obus[data_w*2 +:data_w];
assign c965ibus[temp_w*3 +:temp_w] = v918obus[temp_w*5 +:temp_w];
assign v918ibus[data_w*5 +:data_w] = c965obus[data_w*3 +:data_w];
assign c965ibus[temp_w*4 +:temp_w] = v2117obus[temp_w*1 +:temp_w];
assign v2117ibus[data_w*1 +:data_w] = c965obus[data_w*4 +:data_w];
assign c965ibus[temp_w*5 +:temp_w] = v2213obus[temp_w*0 +:temp_w];
assign v2213ibus[data_w*0 +:data_w] = c965obus[data_w*5 +:data_w];
assign c966ibus[temp_w*0 +:temp_w] = v205obus[temp_w*5 +:temp_w];
assign v205ibus[data_w*5 +:data_w] = c966obus[data_w*0 +:data_w];
assign c966ibus[temp_w*1 +:temp_w] = v359obus[temp_w*2 +:temp_w];
assign v359ibus[data_w*2 +:data_w] = c966obus[data_w*1 +:data_w];
assign c966ibus[temp_w*2 +:temp_w] = v813obus[temp_w*2 +:temp_w];
assign v813ibus[data_w*2 +:data_w] = c966obus[data_w*2 +:data_w];
assign c966ibus[temp_w*3 +:temp_w] = v919obus[temp_w*5 +:temp_w];
assign v919ibus[data_w*5 +:data_w] = c966obus[data_w*3 +:data_w];
assign c966ibus[temp_w*4 +:temp_w] = v2118obus[temp_w*1 +:temp_w];
assign v2118ibus[data_w*1 +:data_w] = c966obus[data_w*4 +:data_w];
assign c966ibus[temp_w*5 +:temp_w] = v2214obus[temp_w*0 +:temp_w];
assign v2214ibus[data_w*0 +:data_w] = c966obus[data_w*5 +:data_w];
assign c967ibus[temp_w*0 +:temp_w] = v206obus[temp_w*5 +:temp_w];
assign v206ibus[data_w*5 +:data_w] = c967obus[data_w*0 +:data_w];
assign c967ibus[temp_w*1 +:temp_w] = v360obus[temp_w*2 +:temp_w];
assign v360ibus[data_w*2 +:data_w] = c967obus[data_w*1 +:data_w];
assign c967ibus[temp_w*2 +:temp_w] = v814obus[temp_w*2 +:temp_w];
assign v814ibus[data_w*2 +:data_w] = c967obus[data_w*2 +:data_w];
assign c967ibus[temp_w*3 +:temp_w] = v920obus[temp_w*5 +:temp_w];
assign v920ibus[data_w*5 +:data_w] = c967obus[data_w*3 +:data_w];
assign c967ibus[temp_w*4 +:temp_w] = v2119obus[temp_w*1 +:temp_w];
assign v2119ibus[data_w*1 +:data_w] = c967obus[data_w*4 +:data_w];
assign c967ibus[temp_w*5 +:temp_w] = v2215obus[temp_w*0 +:temp_w];
assign v2215ibus[data_w*0 +:data_w] = c967obus[data_w*5 +:data_w];
assign c968ibus[temp_w*0 +:temp_w] = v207obus[temp_w*5 +:temp_w];
assign v207ibus[data_w*5 +:data_w] = c968obus[data_w*0 +:data_w];
assign c968ibus[temp_w*1 +:temp_w] = v361obus[temp_w*2 +:temp_w];
assign v361ibus[data_w*2 +:data_w] = c968obus[data_w*1 +:data_w];
assign c968ibus[temp_w*2 +:temp_w] = v815obus[temp_w*2 +:temp_w];
assign v815ibus[data_w*2 +:data_w] = c968obus[data_w*2 +:data_w];
assign c968ibus[temp_w*3 +:temp_w] = v921obus[temp_w*5 +:temp_w];
assign v921ibus[data_w*5 +:data_w] = c968obus[data_w*3 +:data_w];
assign c968ibus[temp_w*4 +:temp_w] = v2120obus[temp_w*1 +:temp_w];
assign v2120ibus[data_w*1 +:data_w] = c968obus[data_w*4 +:data_w];
assign c968ibus[temp_w*5 +:temp_w] = v2216obus[temp_w*0 +:temp_w];
assign v2216ibus[data_w*0 +:data_w] = c968obus[data_w*5 +:data_w];
assign c969ibus[temp_w*0 +:temp_w] = v208obus[temp_w*5 +:temp_w];
assign v208ibus[data_w*5 +:data_w] = c969obus[data_w*0 +:data_w];
assign c969ibus[temp_w*1 +:temp_w] = v362obus[temp_w*2 +:temp_w];
assign v362ibus[data_w*2 +:data_w] = c969obus[data_w*1 +:data_w];
assign c969ibus[temp_w*2 +:temp_w] = v816obus[temp_w*2 +:temp_w];
assign v816ibus[data_w*2 +:data_w] = c969obus[data_w*2 +:data_w];
assign c969ibus[temp_w*3 +:temp_w] = v922obus[temp_w*5 +:temp_w];
assign v922ibus[data_w*5 +:data_w] = c969obus[data_w*3 +:data_w];
assign c969ibus[temp_w*4 +:temp_w] = v2121obus[temp_w*1 +:temp_w];
assign v2121ibus[data_w*1 +:data_w] = c969obus[data_w*4 +:data_w];
assign c969ibus[temp_w*5 +:temp_w] = v2217obus[temp_w*0 +:temp_w];
assign v2217ibus[data_w*0 +:data_w] = c969obus[data_w*5 +:data_w];
assign c970ibus[temp_w*0 +:temp_w] = v209obus[temp_w*5 +:temp_w];
assign v209ibus[data_w*5 +:data_w] = c970obus[data_w*0 +:data_w];
assign c970ibus[temp_w*1 +:temp_w] = v363obus[temp_w*2 +:temp_w];
assign v363ibus[data_w*2 +:data_w] = c970obus[data_w*1 +:data_w];
assign c970ibus[temp_w*2 +:temp_w] = v817obus[temp_w*2 +:temp_w];
assign v817ibus[data_w*2 +:data_w] = c970obus[data_w*2 +:data_w];
assign c970ibus[temp_w*3 +:temp_w] = v923obus[temp_w*5 +:temp_w];
assign v923ibus[data_w*5 +:data_w] = c970obus[data_w*3 +:data_w];
assign c970ibus[temp_w*4 +:temp_w] = v2122obus[temp_w*1 +:temp_w];
assign v2122ibus[data_w*1 +:data_w] = c970obus[data_w*4 +:data_w];
assign c970ibus[temp_w*5 +:temp_w] = v2218obus[temp_w*0 +:temp_w];
assign v2218ibus[data_w*0 +:data_w] = c970obus[data_w*5 +:data_w];
assign c971ibus[temp_w*0 +:temp_w] = v210obus[temp_w*5 +:temp_w];
assign v210ibus[data_w*5 +:data_w] = c971obus[data_w*0 +:data_w];
assign c971ibus[temp_w*1 +:temp_w] = v364obus[temp_w*2 +:temp_w];
assign v364ibus[data_w*2 +:data_w] = c971obus[data_w*1 +:data_w];
assign c971ibus[temp_w*2 +:temp_w] = v818obus[temp_w*2 +:temp_w];
assign v818ibus[data_w*2 +:data_w] = c971obus[data_w*2 +:data_w];
assign c971ibus[temp_w*3 +:temp_w] = v924obus[temp_w*5 +:temp_w];
assign v924ibus[data_w*5 +:data_w] = c971obus[data_w*3 +:data_w];
assign c971ibus[temp_w*4 +:temp_w] = v2123obus[temp_w*1 +:temp_w];
assign v2123ibus[data_w*1 +:data_w] = c971obus[data_w*4 +:data_w];
assign c971ibus[temp_w*5 +:temp_w] = v2219obus[temp_w*0 +:temp_w];
assign v2219ibus[data_w*0 +:data_w] = c971obus[data_w*5 +:data_w];
assign c972ibus[temp_w*0 +:temp_w] = v211obus[temp_w*5 +:temp_w];
assign v211ibus[data_w*5 +:data_w] = c972obus[data_w*0 +:data_w];
assign c972ibus[temp_w*1 +:temp_w] = v365obus[temp_w*2 +:temp_w];
assign v365ibus[data_w*2 +:data_w] = c972obus[data_w*1 +:data_w];
assign c972ibus[temp_w*2 +:temp_w] = v819obus[temp_w*2 +:temp_w];
assign v819ibus[data_w*2 +:data_w] = c972obus[data_w*2 +:data_w];
assign c972ibus[temp_w*3 +:temp_w] = v925obus[temp_w*5 +:temp_w];
assign v925ibus[data_w*5 +:data_w] = c972obus[data_w*3 +:data_w];
assign c972ibus[temp_w*4 +:temp_w] = v2124obus[temp_w*1 +:temp_w];
assign v2124ibus[data_w*1 +:data_w] = c972obus[data_w*4 +:data_w];
assign c972ibus[temp_w*5 +:temp_w] = v2220obus[temp_w*0 +:temp_w];
assign v2220ibus[data_w*0 +:data_w] = c972obus[data_w*5 +:data_w];
assign c973ibus[temp_w*0 +:temp_w] = v212obus[temp_w*5 +:temp_w];
assign v212ibus[data_w*5 +:data_w] = c973obus[data_w*0 +:data_w];
assign c973ibus[temp_w*1 +:temp_w] = v366obus[temp_w*2 +:temp_w];
assign v366ibus[data_w*2 +:data_w] = c973obus[data_w*1 +:data_w];
assign c973ibus[temp_w*2 +:temp_w] = v820obus[temp_w*2 +:temp_w];
assign v820ibus[data_w*2 +:data_w] = c973obus[data_w*2 +:data_w];
assign c973ibus[temp_w*3 +:temp_w] = v926obus[temp_w*5 +:temp_w];
assign v926ibus[data_w*5 +:data_w] = c973obus[data_w*3 +:data_w];
assign c973ibus[temp_w*4 +:temp_w] = v2125obus[temp_w*1 +:temp_w];
assign v2125ibus[data_w*1 +:data_w] = c973obus[data_w*4 +:data_w];
assign c973ibus[temp_w*5 +:temp_w] = v2221obus[temp_w*0 +:temp_w];
assign v2221ibus[data_w*0 +:data_w] = c973obus[data_w*5 +:data_w];
assign c974ibus[temp_w*0 +:temp_w] = v213obus[temp_w*5 +:temp_w];
assign v213ibus[data_w*5 +:data_w] = c974obus[data_w*0 +:data_w];
assign c974ibus[temp_w*1 +:temp_w] = v367obus[temp_w*2 +:temp_w];
assign v367ibus[data_w*2 +:data_w] = c974obus[data_w*1 +:data_w];
assign c974ibus[temp_w*2 +:temp_w] = v821obus[temp_w*2 +:temp_w];
assign v821ibus[data_w*2 +:data_w] = c974obus[data_w*2 +:data_w];
assign c974ibus[temp_w*3 +:temp_w] = v927obus[temp_w*5 +:temp_w];
assign v927ibus[data_w*5 +:data_w] = c974obus[data_w*3 +:data_w];
assign c974ibus[temp_w*4 +:temp_w] = v2126obus[temp_w*1 +:temp_w];
assign v2126ibus[data_w*1 +:data_w] = c974obus[data_w*4 +:data_w];
assign c974ibus[temp_w*5 +:temp_w] = v2222obus[temp_w*0 +:temp_w];
assign v2222ibus[data_w*0 +:data_w] = c974obus[data_w*5 +:data_w];
assign c975ibus[temp_w*0 +:temp_w] = v214obus[temp_w*5 +:temp_w];
assign v214ibus[data_w*5 +:data_w] = c975obus[data_w*0 +:data_w];
assign c975ibus[temp_w*1 +:temp_w] = v368obus[temp_w*2 +:temp_w];
assign v368ibus[data_w*2 +:data_w] = c975obus[data_w*1 +:data_w];
assign c975ibus[temp_w*2 +:temp_w] = v822obus[temp_w*2 +:temp_w];
assign v822ibus[data_w*2 +:data_w] = c975obus[data_w*2 +:data_w];
assign c975ibus[temp_w*3 +:temp_w] = v928obus[temp_w*5 +:temp_w];
assign v928ibus[data_w*5 +:data_w] = c975obus[data_w*3 +:data_w];
assign c975ibus[temp_w*4 +:temp_w] = v2127obus[temp_w*1 +:temp_w];
assign v2127ibus[data_w*1 +:data_w] = c975obus[data_w*4 +:data_w];
assign c975ibus[temp_w*5 +:temp_w] = v2223obus[temp_w*0 +:temp_w];
assign v2223ibus[data_w*0 +:data_w] = c975obus[data_w*5 +:data_w];
assign c976ibus[temp_w*0 +:temp_w] = v215obus[temp_w*5 +:temp_w];
assign v215ibus[data_w*5 +:data_w] = c976obus[data_w*0 +:data_w];
assign c976ibus[temp_w*1 +:temp_w] = v369obus[temp_w*2 +:temp_w];
assign v369ibus[data_w*2 +:data_w] = c976obus[data_w*1 +:data_w];
assign c976ibus[temp_w*2 +:temp_w] = v823obus[temp_w*2 +:temp_w];
assign v823ibus[data_w*2 +:data_w] = c976obus[data_w*2 +:data_w];
assign c976ibus[temp_w*3 +:temp_w] = v929obus[temp_w*5 +:temp_w];
assign v929ibus[data_w*5 +:data_w] = c976obus[data_w*3 +:data_w];
assign c976ibus[temp_w*4 +:temp_w] = v2128obus[temp_w*1 +:temp_w];
assign v2128ibus[data_w*1 +:data_w] = c976obus[data_w*4 +:data_w];
assign c976ibus[temp_w*5 +:temp_w] = v2224obus[temp_w*0 +:temp_w];
assign v2224ibus[data_w*0 +:data_w] = c976obus[data_w*5 +:data_w];
assign c977ibus[temp_w*0 +:temp_w] = v216obus[temp_w*5 +:temp_w];
assign v216ibus[data_w*5 +:data_w] = c977obus[data_w*0 +:data_w];
assign c977ibus[temp_w*1 +:temp_w] = v370obus[temp_w*2 +:temp_w];
assign v370ibus[data_w*2 +:data_w] = c977obus[data_w*1 +:data_w];
assign c977ibus[temp_w*2 +:temp_w] = v824obus[temp_w*2 +:temp_w];
assign v824ibus[data_w*2 +:data_w] = c977obus[data_w*2 +:data_w];
assign c977ibus[temp_w*3 +:temp_w] = v930obus[temp_w*5 +:temp_w];
assign v930ibus[data_w*5 +:data_w] = c977obus[data_w*3 +:data_w];
assign c977ibus[temp_w*4 +:temp_w] = v2129obus[temp_w*1 +:temp_w];
assign v2129ibus[data_w*1 +:data_w] = c977obus[data_w*4 +:data_w];
assign c977ibus[temp_w*5 +:temp_w] = v2225obus[temp_w*0 +:temp_w];
assign v2225ibus[data_w*0 +:data_w] = c977obus[data_w*5 +:data_w];
assign c978ibus[temp_w*0 +:temp_w] = v217obus[temp_w*5 +:temp_w];
assign v217ibus[data_w*5 +:data_w] = c978obus[data_w*0 +:data_w];
assign c978ibus[temp_w*1 +:temp_w] = v371obus[temp_w*2 +:temp_w];
assign v371ibus[data_w*2 +:data_w] = c978obus[data_w*1 +:data_w];
assign c978ibus[temp_w*2 +:temp_w] = v825obus[temp_w*2 +:temp_w];
assign v825ibus[data_w*2 +:data_w] = c978obus[data_w*2 +:data_w];
assign c978ibus[temp_w*3 +:temp_w] = v931obus[temp_w*5 +:temp_w];
assign v931ibus[data_w*5 +:data_w] = c978obus[data_w*3 +:data_w];
assign c978ibus[temp_w*4 +:temp_w] = v2130obus[temp_w*1 +:temp_w];
assign v2130ibus[data_w*1 +:data_w] = c978obus[data_w*4 +:data_w];
assign c978ibus[temp_w*5 +:temp_w] = v2226obus[temp_w*0 +:temp_w];
assign v2226ibus[data_w*0 +:data_w] = c978obus[data_w*5 +:data_w];
assign c979ibus[temp_w*0 +:temp_w] = v218obus[temp_w*5 +:temp_w];
assign v218ibus[data_w*5 +:data_w] = c979obus[data_w*0 +:data_w];
assign c979ibus[temp_w*1 +:temp_w] = v372obus[temp_w*2 +:temp_w];
assign v372ibus[data_w*2 +:data_w] = c979obus[data_w*1 +:data_w];
assign c979ibus[temp_w*2 +:temp_w] = v826obus[temp_w*2 +:temp_w];
assign v826ibus[data_w*2 +:data_w] = c979obus[data_w*2 +:data_w];
assign c979ibus[temp_w*3 +:temp_w] = v932obus[temp_w*5 +:temp_w];
assign v932ibus[data_w*5 +:data_w] = c979obus[data_w*3 +:data_w];
assign c979ibus[temp_w*4 +:temp_w] = v2131obus[temp_w*1 +:temp_w];
assign v2131ibus[data_w*1 +:data_w] = c979obus[data_w*4 +:data_w];
assign c979ibus[temp_w*5 +:temp_w] = v2227obus[temp_w*0 +:temp_w];
assign v2227ibus[data_w*0 +:data_w] = c979obus[data_w*5 +:data_w];
assign c980ibus[temp_w*0 +:temp_w] = v219obus[temp_w*5 +:temp_w];
assign v219ibus[data_w*5 +:data_w] = c980obus[data_w*0 +:data_w];
assign c980ibus[temp_w*1 +:temp_w] = v373obus[temp_w*2 +:temp_w];
assign v373ibus[data_w*2 +:data_w] = c980obus[data_w*1 +:data_w];
assign c980ibus[temp_w*2 +:temp_w] = v827obus[temp_w*2 +:temp_w];
assign v827ibus[data_w*2 +:data_w] = c980obus[data_w*2 +:data_w];
assign c980ibus[temp_w*3 +:temp_w] = v933obus[temp_w*5 +:temp_w];
assign v933ibus[data_w*5 +:data_w] = c980obus[data_w*3 +:data_w];
assign c980ibus[temp_w*4 +:temp_w] = v2132obus[temp_w*1 +:temp_w];
assign v2132ibus[data_w*1 +:data_w] = c980obus[data_w*4 +:data_w];
assign c980ibus[temp_w*5 +:temp_w] = v2228obus[temp_w*0 +:temp_w];
assign v2228ibus[data_w*0 +:data_w] = c980obus[data_w*5 +:data_w];
assign c981ibus[temp_w*0 +:temp_w] = v220obus[temp_w*5 +:temp_w];
assign v220ibus[data_w*5 +:data_w] = c981obus[data_w*0 +:data_w];
assign c981ibus[temp_w*1 +:temp_w] = v374obus[temp_w*2 +:temp_w];
assign v374ibus[data_w*2 +:data_w] = c981obus[data_w*1 +:data_w];
assign c981ibus[temp_w*2 +:temp_w] = v828obus[temp_w*2 +:temp_w];
assign v828ibus[data_w*2 +:data_w] = c981obus[data_w*2 +:data_w];
assign c981ibus[temp_w*3 +:temp_w] = v934obus[temp_w*5 +:temp_w];
assign v934ibus[data_w*5 +:data_w] = c981obus[data_w*3 +:data_w];
assign c981ibus[temp_w*4 +:temp_w] = v2133obus[temp_w*1 +:temp_w];
assign v2133ibus[data_w*1 +:data_w] = c981obus[data_w*4 +:data_w];
assign c981ibus[temp_w*5 +:temp_w] = v2229obus[temp_w*0 +:temp_w];
assign v2229ibus[data_w*0 +:data_w] = c981obus[data_w*5 +:data_w];
assign c982ibus[temp_w*0 +:temp_w] = v221obus[temp_w*5 +:temp_w];
assign v221ibus[data_w*5 +:data_w] = c982obus[data_w*0 +:data_w];
assign c982ibus[temp_w*1 +:temp_w] = v375obus[temp_w*2 +:temp_w];
assign v375ibus[data_w*2 +:data_w] = c982obus[data_w*1 +:data_w];
assign c982ibus[temp_w*2 +:temp_w] = v829obus[temp_w*2 +:temp_w];
assign v829ibus[data_w*2 +:data_w] = c982obus[data_w*2 +:data_w];
assign c982ibus[temp_w*3 +:temp_w] = v935obus[temp_w*5 +:temp_w];
assign v935ibus[data_w*5 +:data_w] = c982obus[data_w*3 +:data_w];
assign c982ibus[temp_w*4 +:temp_w] = v2134obus[temp_w*1 +:temp_w];
assign v2134ibus[data_w*1 +:data_w] = c982obus[data_w*4 +:data_w];
assign c982ibus[temp_w*5 +:temp_w] = v2230obus[temp_w*0 +:temp_w];
assign v2230ibus[data_w*0 +:data_w] = c982obus[data_w*5 +:data_w];
assign c983ibus[temp_w*0 +:temp_w] = v222obus[temp_w*5 +:temp_w];
assign v222ibus[data_w*5 +:data_w] = c983obus[data_w*0 +:data_w];
assign c983ibus[temp_w*1 +:temp_w] = v376obus[temp_w*2 +:temp_w];
assign v376ibus[data_w*2 +:data_w] = c983obus[data_w*1 +:data_w];
assign c983ibus[temp_w*2 +:temp_w] = v830obus[temp_w*2 +:temp_w];
assign v830ibus[data_w*2 +:data_w] = c983obus[data_w*2 +:data_w];
assign c983ibus[temp_w*3 +:temp_w] = v936obus[temp_w*5 +:temp_w];
assign v936ibus[data_w*5 +:data_w] = c983obus[data_w*3 +:data_w];
assign c983ibus[temp_w*4 +:temp_w] = v2135obus[temp_w*1 +:temp_w];
assign v2135ibus[data_w*1 +:data_w] = c983obus[data_w*4 +:data_w];
assign c983ibus[temp_w*5 +:temp_w] = v2231obus[temp_w*0 +:temp_w];
assign v2231ibus[data_w*0 +:data_w] = c983obus[data_w*5 +:data_w];
assign c984ibus[temp_w*0 +:temp_w] = v223obus[temp_w*5 +:temp_w];
assign v223ibus[data_w*5 +:data_w] = c984obus[data_w*0 +:data_w];
assign c984ibus[temp_w*1 +:temp_w] = v377obus[temp_w*2 +:temp_w];
assign v377ibus[data_w*2 +:data_w] = c984obus[data_w*1 +:data_w];
assign c984ibus[temp_w*2 +:temp_w] = v831obus[temp_w*2 +:temp_w];
assign v831ibus[data_w*2 +:data_w] = c984obus[data_w*2 +:data_w];
assign c984ibus[temp_w*3 +:temp_w] = v937obus[temp_w*5 +:temp_w];
assign v937ibus[data_w*5 +:data_w] = c984obus[data_w*3 +:data_w];
assign c984ibus[temp_w*4 +:temp_w] = v2136obus[temp_w*1 +:temp_w];
assign v2136ibus[data_w*1 +:data_w] = c984obus[data_w*4 +:data_w];
assign c984ibus[temp_w*5 +:temp_w] = v2232obus[temp_w*0 +:temp_w];
assign v2232ibus[data_w*0 +:data_w] = c984obus[data_w*5 +:data_w];
assign c985ibus[temp_w*0 +:temp_w] = v224obus[temp_w*5 +:temp_w];
assign v224ibus[data_w*5 +:data_w] = c985obus[data_w*0 +:data_w];
assign c985ibus[temp_w*1 +:temp_w] = v378obus[temp_w*2 +:temp_w];
assign v378ibus[data_w*2 +:data_w] = c985obus[data_w*1 +:data_w];
assign c985ibus[temp_w*2 +:temp_w] = v832obus[temp_w*2 +:temp_w];
assign v832ibus[data_w*2 +:data_w] = c985obus[data_w*2 +:data_w];
assign c985ibus[temp_w*3 +:temp_w] = v938obus[temp_w*5 +:temp_w];
assign v938ibus[data_w*5 +:data_w] = c985obus[data_w*3 +:data_w];
assign c985ibus[temp_w*4 +:temp_w] = v2137obus[temp_w*1 +:temp_w];
assign v2137ibus[data_w*1 +:data_w] = c985obus[data_w*4 +:data_w];
assign c985ibus[temp_w*5 +:temp_w] = v2233obus[temp_w*0 +:temp_w];
assign v2233ibus[data_w*0 +:data_w] = c985obus[data_w*5 +:data_w];
assign c986ibus[temp_w*0 +:temp_w] = v225obus[temp_w*5 +:temp_w];
assign v225ibus[data_w*5 +:data_w] = c986obus[data_w*0 +:data_w];
assign c986ibus[temp_w*1 +:temp_w] = v379obus[temp_w*2 +:temp_w];
assign v379ibus[data_w*2 +:data_w] = c986obus[data_w*1 +:data_w];
assign c986ibus[temp_w*2 +:temp_w] = v833obus[temp_w*2 +:temp_w];
assign v833ibus[data_w*2 +:data_w] = c986obus[data_w*2 +:data_w];
assign c986ibus[temp_w*3 +:temp_w] = v939obus[temp_w*5 +:temp_w];
assign v939ibus[data_w*5 +:data_w] = c986obus[data_w*3 +:data_w];
assign c986ibus[temp_w*4 +:temp_w] = v2138obus[temp_w*1 +:temp_w];
assign v2138ibus[data_w*1 +:data_w] = c986obus[data_w*4 +:data_w];
assign c986ibus[temp_w*5 +:temp_w] = v2234obus[temp_w*0 +:temp_w];
assign v2234ibus[data_w*0 +:data_w] = c986obus[data_w*5 +:data_w];
assign c987ibus[temp_w*0 +:temp_w] = v226obus[temp_w*5 +:temp_w];
assign v226ibus[data_w*5 +:data_w] = c987obus[data_w*0 +:data_w];
assign c987ibus[temp_w*1 +:temp_w] = v380obus[temp_w*2 +:temp_w];
assign v380ibus[data_w*2 +:data_w] = c987obus[data_w*1 +:data_w];
assign c987ibus[temp_w*2 +:temp_w] = v834obus[temp_w*2 +:temp_w];
assign v834ibus[data_w*2 +:data_w] = c987obus[data_w*2 +:data_w];
assign c987ibus[temp_w*3 +:temp_w] = v940obus[temp_w*5 +:temp_w];
assign v940ibus[data_w*5 +:data_w] = c987obus[data_w*3 +:data_w];
assign c987ibus[temp_w*4 +:temp_w] = v2139obus[temp_w*1 +:temp_w];
assign v2139ibus[data_w*1 +:data_w] = c987obus[data_w*4 +:data_w];
assign c987ibus[temp_w*5 +:temp_w] = v2235obus[temp_w*0 +:temp_w];
assign v2235ibus[data_w*0 +:data_w] = c987obus[data_w*5 +:data_w];
assign c988ibus[temp_w*0 +:temp_w] = v227obus[temp_w*5 +:temp_w];
assign v227ibus[data_w*5 +:data_w] = c988obus[data_w*0 +:data_w];
assign c988ibus[temp_w*1 +:temp_w] = v381obus[temp_w*2 +:temp_w];
assign v381ibus[data_w*2 +:data_w] = c988obus[data_w*1 +:data_w];
assign c988ibus[temp_w*2 +:temp_w] = v835obus[temp_w*2 +:temp_w];
assign v835ibus[data_w*2 +:data_w] = c988obus[data_w*2 +:data_w];
assign c988ibus[temp_w*3 +:temp_w] = v941obus[temp_w*5 +:temp_w];
assign v941ibus[data_w*5 +:data_w] = c988obus[data_w*3 +:data_w];
assign c988ibus[temp_w*4 +:temp_w] = v2140obus[temp_w*1 +:temp_w];
assign v2140ibus[data_w*1 +:data_w] = c988obus[data_w*4 +:data_w];
assign c988ibus[temp_w*5 +:temp_w] = v2236obus[temp_w*0 +:temp_w];
assign v2236ibus[data_w*0 +:data_w] = c988obus[data_w*5 +:data_w];
assign c989ibus[temp_w*0 +:temp_w] = v228obus[temp_w*5 +:temp_w];
assign v228ibus[data_w*5 +:data_w] = c989obus[data_w*0 +:data_w];
assign c989ibus[temp_w*1 +:temp_w] = v382obus[temp_w*2 +:temp_w];
assign v382ibus[data_w*2 +:data_w] = c989obus[data_w*1 +:data_w];
assign c989ibus[temp_w*2 +:temp_w] = v836obus[temp_w*2 +:temp_w];
assign v836ibus[data_w*2 +:data_w] = c989obus[data_w*2 +:data_w];
assign c989ibus[temp_w*3 +:temp_w] = v942obus[temp_w*5 +:temp_w];
assign v942ibus[data_w*5 +:data_w] = c989obus[data_w*3 +:data_w];
assign c989ibus[temp_w*4 +:temp_w] = v2141obus[temp_w*1 +:temp_w];
assign v2141ibus[data_w*1 +:data_w] = c989obus[data_w*4 +:data_w];
assign c989ibus[temp_w*5 +:temp_w] = v2237obus[temp_w*0 +:temp_w];
assign v2237ibus[data_w*0 +:data_w] = c989obus[data_w*5 +:data_w];
assign c990ibus[temp_w*0 +:temp_w] = v229obus[temp_w*5 +:temp_w];
assign v229ibus[data_w*5 +:data_w] = c990obus[data_w*0 +:data_w];
assign c990ibus[temp_w*1 +:temp_w] = v383obus[temp_w*2 +:temp_w];
assign v383ibus[data_w*2 +:data_w] = c990obus[data_w*1 +:data_w];
assign c990ibus[temp_w*2 +:temp_w] = v837obus[temp_w*2 +:temp_w];
assign v837ibus[data_w*2 +:data_w] = c990obus[data_w*2 +:data_w];
assign c990ibus[temp_w*3 +:temp_w] = v943obus[temp_w*5 +:temp_w];
assign v943ibus[data_w*5 +:data_w] = c990obus[data_w*3 +:data_w];
assign c990ibus[temp_w*4 +:temp_w] = v2142obus[temp_w*1 +:temp_w];
assign v2142ibus[data_w*1 +:data_w] = c990obus[data_w*4 +:data_w];
assign c990ibus[temp_w*5 +:temp_w] = v2238obus[temp_w*0 +:temp_w];
assign v2238ibus[data_w*0 +:data_w] = c990obus[data_w*5 +:data_w];
assign c991ibus[temp_w*0 +:temp_w] = v230obus[temp_w*5 +:temp_w];
assign v230ibus[data_w*5 +:data_w] = c991obus[data_w*0 +:data_w];
assign c991ibus[temp_w*1 +:temp_w] = v288obus[temp_w*2 +:temp_w];
assign v288ibus[data_w*2 +:data_w] = c991obus[data_w*1 +:data_w];
assign c991ibus[temp_w*2 +:temp_w] = v838obus[temp_w*2 +:temp_w];
assign v838ibus[data_w*2 +:data_w] = c991obus[data_w*2 +:data_w];
assign c991ibus[temp_w*3 +:temp_w] = v944obus[temp_w*5 +:temp_w];
assign v944ibus[data_w*5 +:data_w] = c991obus[data_w*3 +:data_w];
assign c991ibus[temp_w*4 +:temp_w] = v2143obus[temp_w*1 +:temp_w];
assign v2143ibus[data_w*1 +:data_w] = c991obus[data_w*4 +:data_w];
assign c991ibus[temp_w*5 +:temp_w] = v2239obus[temp_w*0 +:temp_w];
assign v2239ibus[data_w*0 +:data_w] = c991obus[data_w*5 +:data_w];
assign c992ibus[temp_w*0 +:temp_w] = v231obus[temp_w*5 +:temp_w];
assign v231ibus[data_w*5 +:data_w] = c992obus[data_w*0 +:data_w];
assign c992ibus[temp_w*1 +:temp_w] = v289obus[temp_w*2 +:temp_w];
assign v289ibus[data_w*2 +:data_w] = c992obus[data_w*1 +:data_w];
assign c992ibus[temp_w*2 +:temp_w] = v839obus[temp_w*2 +:temp_w];
assign v839ibus[data_w*2 +:data_w] = c992obus[data_w*2 +:data_w];
assign c992ibus[temp_w*3 +:temp_w] = v945obus[temp_w*5 +:temp_w];
assign v945ibus[data_w*5 +:data_w] = c992obus[data_w*3 +:data_w];
assign c992ibus[temp_w*4 +:temp_w] = v2144obus[temp_w*1 +:temp_w];
assign v2144ibus[data_w*1 +:data_w] = c992obus[data_w*4 +:data_w];
assign c992ibus[temp_w*5 +:temp_w] = v2240obus[temp_w*0 +:temp_w];
assign v2240ibus[data_w*0 +:data_w] = c992obus[data_w*5 +:data_w];
assign c993ibus[temp_w*0 +:temp_w] = v232obus[temp_w*5 +:temp_w];
assign v232ibus[data_w*5 +:data_w] = c993obus[data_w*0 +:data_w];
assign c993ibus[temp_w*1 +:temp_w] = v290obus[temp_w*2 +:temp_w];
assign v290ibus[data_w*2 +:data_w] = c993obus[data_w*1 +:data_w];
assign c993ibus[temp_w*2 +:temp_w] = v840obus[temp_w*2 +:temp_w];
assign v840ibus[data_w*2 +:data_w] = c993obus[data_w*2 +:data_w];
assign c993ibus[temp_w*3 +:temp_w] = v946obus[temp_w*5 +:temp_w];
assign v946ibus[data_w*5 +:data_w] = c993obus[data_w*3 +:data_w];
assign c993ibus[temp_w*4 +:temp_w] = v2145obus[temp_w*1 +:temp_w];
assign v2145ibus[data_w*1 +:data_w] = c993obus[data_w*4 +:data_w];
assign c993ibus[temp_w*5 +:temp_w] = v2241obus[temp_w*0 +:temp_w];
assign v2241ibus[data_w*0 +:data_w] = c993obus[data_w*5 +:data_w];
assign c994ibus[temp_w*0 +:temp_w] = v233obus[temp_w*5 +:temp_w];
assign v233ibus[data_w*5 +:data_w] = c994obus[data_w*0 +:data_w];
assign c994ibus[temp_w*1 +:temp_w] = v291obus[temp_w*2 +:temp_w];
assign v291ibus[data_w*2 +:data_w] = c994obus[data_w*1 +:data_w];
assign c994ibus[temp_w*2 +:temp_w] = v841obus[temp_w*2 +:temp_w];
assign v841ibus[data_w*2 +:data_w] = c994obus[data_w*2 +:data_w];
assign c994ibus[temp_w*3 +:temp_w] = v947obus[temp_w*5 +:temp_w];
assign v947ibus[data_w*5 +:data_w] = c994obus[data_w*3 +:data_w];
assign c994ibus[temp_w*4 +:temp_w] = v2146obus[temp_w*1 +:temp_w];
assign v2146ibus[data_w*1 +:data_w] = c994obus[data_w*4 +:data_w];
assign c994ibus[temp_w*5 +:temp_w] = v2242obus[temp_w*0 +:temp_w];
assign v2242ibus[data_w*0 +:data_w] = c994obus[data_w*5 +:data_w];
assign c995ibus[temp_w*0 +:temp_w] = v234obus[temp_w*5 +:temp_w];
assign v234ibus[data_w*5 +:data_w] = c995obus[data_w*0 +:data_w];
assign c995ibus[temp_w*1 +:temp_w] = v292obus[temp_w*2 +:temp_w];
assign v292ibus[data_w*2 +:data_w] = c995obus[data_w*1 +:data_w];
assign c995ibus[temp_w*2 +:temp_w] = v842obus[temp_w*2 +:temp_w];
assign v842ibus[data_w*2 +:data_w] = c995obus[data_w*2 +:data_w];
assign c995ibus[temp_w*3 +:temp_w] = v948obus[temp_w*5 +:temp_w];
assign v948ibus[data_w*5 +:data_w] = c995obus[data_w*3 +:data_w];
assign c995ibus[temp_w*4 +:temp_w] = v2147obus[temp_w*1 +:temp_w];
assign v2147ibus[data_w*1 +:data_w] = c995obus[data_w*4 +:data_w];
assign c995ibus[temp_w*5 +:temp_w] = v2243obus[temp_w*0 +:temp_w];
assign v2243ibus[data_w*0 +:data_w] = c995obus[data_w*5 +:data_w];
assign c996ibus[temp_w*0 +:temp_w] = v235obus[temp_w*5 +:temp_w];
assign v235ibus[data_w*5 +:data_w] = c996obus[data_w*0 +:data_w];
assign c996ibus[temp_w*1 +:temp_w] = v293obus[temp_w*2 +:temp_w];
assign v293ibus[data_w*2 +:data_w] = c996obus[data_w*1 +:data_w];
assign c996ibus[temp_w*2 +:temp_w] = v843obus[temp_w*2 +:temp_w];
assign v843ibus[data_w*2 +:data_w] = c996obus[data_w*2 +:data_w];
assign c996ibus[temp_w*3 +:temp_w] = v949obus[temp_w*5 +:temp_w];
assign v949ibus[data_w*5 +:data_w] = c996obus[data_w*3 +:data_w];
assign c996ibus[temp_w*4 +:temp_w] = v2148obus[temp_w*1 +:temp_w];
assign v2148ibus[data_w*1 +:data_w] = c996obus[data_w*4 +:data_w];
assign c996ibus[temp_w*5 +:temp_w] = v2244obus[temp_w*0 +:temp_w];
assign v2244ibus[data_w*0 +:data_w] = c996obus[data_w*5 +:data_w];
assign c997ibus[temp_w*0 +:temp_w] = v236obus[temp_w*5 +:temp_w];
assign v236ibus[data_w*5 +:data_w] = c997obus[data_w*0 +:data_w];
assign c997ibus[temp_w*1 +:temp_w] = v294obus[temp_w*2 +:temp_w];
assign v294ibus[data_w*2 +:data_w] = c997obus[data_w*1 +:data_w];
assign c997ibus[temp_w*2 +:temp_w] = v844obus[temp_w*2 +:temp_w];
assign v844ibus[data_w*2 +:data_w] = c997obus[data_w*2 +:data_w];
assign c997ibus[temp_w*3 +:temp_w] = v950obus[temp_w*5 +:temp_w];
assign v950ibus[data_w*5 +:data_w] = c997obus[data_w*3 +:data_w];
assign c997ibus[temp_w*4 +:temp_w] = v2149obus[temp_w*1 +:temp_w];
assign v2149ibus[data_w*1 +:data_w] = c997obus[data_w*4 +:data_w];
assign c997ibus[temp_w*5 +:temp_w] = v2245obus[temp_w*0 +:temp_w];
assign v2245ibus[data_w*0 +:data_w] = c997obus[data_w*5 +:data_w];
assign c998ibus[temp_w*0 +:temp_w] = v237obus[temp_w*5 +:temp_w];
assign v237ibus[data_w*5 +:data_w] = c998obus[data_w*0 +:data_w];
assign c998ibus[temp_w*1 +:temp_w] = v295obus[temp_w*2 +:temp_w];
assign v295ibus[data_w*2 +:data_w] = c998obus[data_w*1 +:data_w];
assign c998ibus[temp_w*2 +:temp_w] = v845obus[temp_w*2 +:temp_w];
assign v845ibus[data_w*2 +:data_w] = c998obus[data_w*2 +:data_w];
assign c998ibus[temp_w*3 +:temp_w] = v951obus[temp_w*5 +:temp_w];
assign v951ibus[data_w*5 +:data_w] = c998obus[data_w*3 +:data_w];
assign c998ibus[temp_w*4 +:temp_w] = v2150obus[temp_w*1 +:temp_w];
assign v2150ibus[data_w*1 +:data_w] = c998obus[data_w*4 +:data_w];
assign c998ibus[temp_w*5 +:temp_w] = v2246obus[temp_w*0 +:temp_w];
assign v2246ibus[data_w*0 +:data_w] = c998obus[data_w*5 +:data_w];
assign c999ibus[temp_w*0 +:temp_w] = v238obus[temp_w*5 +:temp_w];
assign v238ibus[data_w*5 +:data_w] = c999obus[data_w*0 +:data_w];
assign c999ibus[temp_w*1 +:temp_w] = v296obus[temp_w*2 +:temp_w];
assign v296ibus[data_w*2 +:data_w] = c999obus[data_w*1 +:data_w];
assign c999ibus[temp_w*2 +:temp_w] = v846obus[temp_w*2 +:temp_w];
assign v846ibus[data_w*2 +:data_w] = c999obus[data_w*2 +:data_w];
assign c999ibus[temp_w*3 +:temp_w] = v952obus[temp_w*5 +:temp_w];
assign v952ibus[data_w*5 +:data_w] = c999obus[data_w*3 +:data_w];
assign c999ibus[temp_w*4 +:temp_w] = v2151obus[temp_w*1 +:temp_w];
assign v2151ibus[data_w*1 +:data_w] = c999obus[data_w*4 +:data_w];
assign c999ibus[temp_w*5 +:temp_w] = v2247obus[temp_w*0 +:temp_w];
assign v2247ibus[data_w*0 +:data_w] = c999obus[data_w*5 +:data_w];
assign c1000ibus[temp_w*0 +:temp_w] = v239obus[temp_w*5 +:temp_w];
assign v239ibus[data_w*5 +:data_w] = c1000obus[data_w*0 +:data_w];
assign c1000ibus[temp_w*1 +:temp_w] = v297obus[temp_w*2 +:temp_w];
assign v297ibus[data_w*2 +:data_w] = c1000obus[data_w*1 +:data_w];
assign c1000ibus[temp_w*2 +:temp_w] = v847obus[temp_w*2 +:temp_w];
assign v847ibus[data_w*2 +:data_w] = c1000obus[data_w*2 +:data_w];
assign c1000ibus[temp_w*3 +:temp_w] = v953obus[temp_w*5 +:temp_w];
assign v953ibus[data_w*5 +:data_w] = c1000obus[data_w*3 +:data_w];
assign c1000ibus[temp_w*4 +:temp_w] = v2152obus[temp_w*1 +:temp_w];
assign v2152ibus[data_w*1 +:data_w] = c1000obus[data_w*4 +:data_w];
assign c1000ibus[temp_w*5 +:temp_w] = v2248obus[temp_w*0 +:temp_w];
assign v2248ibus[data_w*0 +:data_w] = c1000obus[data_w*5 +:data_w];
assign c1001ibus[temp_w*0 +:temp_w] = v240obus[temp_w*5 +:temp_w];
assign v240ibus[data_w*5 +:data_w] = c1001obus[data_w*0 +:data_w];
assign c1001ibus[temp_w*1 +:temp_w] = v298obus[temp_w*2 +:temp_w];
assign v298ibus[data_w*2 +:data_w] = c1001obus[data_w*1 +:data_w];
assign c1001ibus[temp_w*2 +:temp_w] = v848obus[temp_w*2 +:temp_w];
assign v848ibus[data_w*2 +:data_w] = c1001obus[data_w*2 +:data_w];
assign c1001ibus[temp_w*3 +:temp_w] = v954obus[temp_w*5 +:temp_w];
assign v954ibus[data_w*5 +:data_w] = c1001obus[data_w*3 +:data_w];
assign c1001ibus[temp_w*4 +:temp_w] = v2153obus[temp_w*1 +:temp_w];
assign v2153ibus[data_w*1 +:data_w] = c1001obus[data_w*4 +:data_w];
assign c1001ibus[temp_w*5 +:temp_w] = v2249obus[temp_w*0 +:temp_w];
assign v2249ibus[data_w*0 +:data_w] = c1001obus[data_w*5 +:data_w];
assign c1002ibus[temp_w*0 +:temp_w] = v241obus[temp_w*5 +:temp_w];
assign v241ibus[data_w*5 +:data_w] = c1002obus[data_w*0 +:data_w];
assign c1002ibus[temp_w*1 +:temp_w] = v299obus[temp_w*2 +:temp_w];
assign v299ibus[data_w*2 +:data_w] = c1002obus[data_w*1 +:data_w];
assign c1002ibus[temp_w*2 +:temp_w] = v849obus[temp_w*2 +:temp_w];
assign v849ibus[data_w*2 +:data_w] = c1002obus[data_w*2 +:data_w];
assign c1002ibus[temp_w*3 +:temp_w] = v955obus[temp_w*5 +:temp_w];
assign v955ibus[data_w*5 +:data_w] = c1002obus[data_w*3 +:data_w];
assign c1002ibus[temp_w*4 +:temp_w] = v2154obus[temp_w*1 +:temp_w];
assign v2154ibus[data_w*1 +:data_w] = c1002obus[data_w*4 +:data_w];
assign c1002ibus[temp_w*5 +:temp_w] = v2250obus[temp_w*0 +:temp_w];
assign v2250ibus[data_w*0 +:data_w] = c1002obus[data_w*5 +:data_w];
assign c1003ibus[temp_w*0 +:temp_w] = v242obus[temp_w*5 +:temp_w];
assign v242ibus[data_w*5 +:data_w] = c1003obus[data_w*0 +:data_w];
assign c1003ibus[temp_w*1 +:temp_w] = v300obus[temp_w*2 +:temp_w];
assign v300ibus[data_w*2 +:data_w] = c1003obus[data_w*1 +:data_w];
assign c1003ibus[temp_w*2 +:temp_w] = v850obus[temp_w*2 +:temp_w];
assign v850ibus[data_w*2 +:data_w] = c1003obus[data_w*2 +:data_w];
assign c1003ibus[temp_w*3 +:temp_w] = v956obus[temp_w*5 +:temp_w];
assign v956ibus[data_w*5 +:data_w] = c1003obus[data_w*3 +:data_w];
assign c1003ibus[temp_w*4 +:temp_w] = v2155obus[temp_w*1 +:temp_w];
assign v2155ibus[data_w*1 +:data_w] = c1003obus[data_w*4 +:data_w];
assign c1003ibus[temp_w*5 +:temp_w] = v2251obus[temp_w*0 +:temp_w];
assign v2251ibus[data_w*0 +:data_w] = c1003obus[data_w*5 +:data_w];
assign c1004ibus[temp_w*0 +:temp_w] = v243obus[temp_w*5 +:temp_w];
assign v243ibus[data_w*5 +:data_w] = c1004obus[data_w*0 +:data_w];
assign c1004ibus[temp_w*1 +:temp_w] = v301obus[temp_w*2 +:temp_w];
assign v301ibus[data_w*2 +:data_w] = c1004obus[data_w*1 +:data_w];
assign c1004ibus[temp_w*2 +:temp_w] = v851obus[temp_w*2 +:temp_w];
assign v851ibus[data_w*2 +:data_w] = c1004obus[data_w*2 +:data_w];
assign c1004ibus[temp_w*3 +:temp_w] = v957obus[temp_w*5 +:temp_w];
assign v957ibus[data_w*5 +:data_w] = c1004obus[data_w*3 +:data_w];
assign c1004ibus[temp_w*4 +:temp_w] = v2156obus[temp_w*1 +:temp_w];
assign v2156ibus[data_w*1 +:data_w] = c1004obus[data_w*4 +:data_w];
assign c1004ibus[temp_w*5 +:temp_w] = v2252obus[temp_w*0 +:temp_w];
assign v2252ibus[data_w*0 +:data_w] = c1004obus[data_w*5 +:data_w];
assign c1005ibus[temp_w*0 +:temp_w] = v244obus[temp_w*5 +:temp_w];
assign v244ibus[data_w*5 +:data_w] = c1005obus[data_w*0 +:data_w];
assign c1005ibus[temp_w*1 +:temp_w] = v302obus[temp_w*2 +:temp_w];
assign v302ibus[data_w*2 +:data_w] = c1005obus[data_w*1 +:data_w];
assign c1005ibus[temp_w*2 +:temp_w] = v852obus[temp_w*2 +:temp_w];
assign v852ibus[data_w*2 +:data_w] = c1005obus[data_w*2 +:data_w];
assign c1005ibus[temp_w*3 +:temp_w] = v958obus[temp_w*5 +:temp_w];
assign v958ibus[data_w*5 +:data_w] = c1005obus[data_w*3 +:data_w];
assign c1005ibus[temp_w*4 +:temp_w] = v2157obus[temp_w*1 +:temp_w];
assign v2157ibus[data_w*1 +:data_w] = c1005obus[data_w*4 +:data_w];
assign c1005ibus[temp_w*5 +:temp_w] = v2253obus[temp_w*0 +:temp_w];
assign v2253ibus[data_w*0 +:data_w] = c1005obus[data_w*5 +:data_w];
assign c1006ibus[temp_w*0 +:temp_w] = v245obus[temp_w*5 +:temp_w];
assign v245ibus[data_w*5 +:data_w] = c1006obus[data_w*0 +:data_w];
assign c1006ibus[temp_w*1 +:temp_w] = v303obus[temp_w*2 +:temp_w];
assign v303ibus[data_w*2 +:data_w] = c1006obus[data_w*1 +:data_w];
assign c1006ibus[temp_w*2 +:temp_w] = v853obus[temp_w*2 +:temp_w];
assign v853ibus[data_w*2 +:data_w] = c1006obus[data_w*2 +:data_w];
assign c1006ibus[temp_w*3 +:temp_w] = v959obus[temp_w*5 +:temp_w];
assign v959ibus[data_w*5 +:data_w] = c1006obus[data_w*3 +:data_w];
assign c1006ibus[temp_w*4 +:temp_w] = v2158obus[temp_w*1 +:temp_w];
assign v2158ibus[data_w*1 +:data_w] = c1006obus[data_w*4 +:data_w];
assign c1006ibus[temp_w*5 +:temp_w] = v2254obus[temp_w*0 +:temp_w];
assign v2254ibus[data_w*0 +:data_w] = c1006obus[data_w*5 +:data_w];
assign c1007ibus[temp_w*0 +:temp_w] = v246obus[temp_w*5 +:temp_w];
assign v246ibus[data_w*5 +:data_w] = c1007obus[data_w*0 +:data_w];
assign c1007ibus[temp_w*1 +:temp_w] = v304obus[temp_w*2 +:temp_w];
assign v304ibus[data_w*2 +:data_w] = c1007obus[data_w*1 +:data_w];
assign c1007ibus[temp_w*2 +:temp_w] = v854obus[temp_w*2 +:temp_w];
assign v854ibus[data_w*2 +:data_w] = c1007obus[data_w*2 +:data_w];
assign c1007ibus[temp_w*3 +:temp_w] = v864obus[temp_w*5 +:temp_w];
assign v864ibus[data_w*5 +:data_w] = c1007obus[data_w*3 +:data_w];
assign c1007ibus[temp_w*4 +:temp_w] = v2159obus[temp_w*1 +:temp_w];
assign v2159ibus[data_w*1 +:data_w] = c1007obus[data_w*4 +:data_w];
assign c1007ibus[temp_w*5 +:temp_w] = v2255obus[temp_w*0 +:temp_w];
assign v2255ibus[data_w*0 +:data_w] = c1007obus[data_w*5 +:data_w];
assign c1008ibus[temp_w*0 +:temp_w] = v247obus[temp_w*5 +:temp_w];
assign v247ibus[data_w*5 +:data_w] = c1008obus[data_w*0 +:data_w];
assign c1008ibus[temp_w*1 +:temp_w] = v305obus[temp_w*2 +:temp_w];
assign v305ibus[data_w*2 +:data_w] = c1008obus[data_w*1 +:data_w];
assign c1008ibus[temp_w*2 +:temp_w] = v855obus[temp_w*2 +:temp_w];
assign v855ibus[data_w*2 +:data_w] = c1008obus[data_w*2 +:data_w];
assign c1008ibus[temp_w*3 +:temp_w] = v865obus[temp_w*5 +:temp_w];
assign v865ibus[data_w*5 +:data_w] = c1008obus[data_w*3 +:data_w];
assign c1008ibus[temp_w*4 +:temp_w] = v2160obus[temp_w*1 +:temp_w];
assign v2160ibus[data_w*1 +:data_w] = c1008obus[data_w*4 +:data_w];
assign c1008ibus[temp_w*5 +:temp_w] = v2256obus[temp_w*0 +:temp_w];
assign v2256ibus[data_w*0 +:data_w] = c1008obus[data_w*5 +:data_w];
assign c1009ibus[temp_w*0 +:temp_w] = v248obus[temp_w*5 +:temp_w];
assign v248ibus[data_w*5 +:data_w] = c1009obus[data_w*0 +:data_w];
assign c1009ibus[temp_w*1 +:temp_w] = v306obus[temp_w*2 +:temp_w];
assign v306ibus[data_w*2 +:data_w] = c1009obus[data_w*1 +:data_w];
assign c1009ibus[temp_w*2 +:temp_w] = v856obus[temp_w*2 +:temp_w];
assign v856ibus[data_w*2 +:data_w] = c1009obus[data_w*2 +:data_w];
assign c1009ibus[temp_w*3 +:temp_w] = v866obus[temp_w*5 +:temp_w];
assign v866ibus[data_w*5 +:data_w] = c1009obus[data_w*3 +:data_w];
assign c1009ibus[temp_w*4 +:temp_w] = v2161obus[temp_w*1 +:temp_w];
assign v2161ibus[data_w*1 +:data_w] = c1009obus[data_w*4 +:data_w];
assign c1009ibus[temp_w*5 +:temp_w] = v2257obus[temp_w*0 +:temp_w];
assign v2257ibus[data_w*0 +:data_w] = c1009obus[data_w*5 +:data_w];
assign c1010ibus[temp_w*0 +:temp_w] = v249obus[temp_w*5 +:temp_w];
assign v249ibus[data_w*5 +:data_w] = c1010obus[data_w*0 +:data_w];
assign c1010ibus[temp_w*1 +:temp_w] = v307obus[temp_w*2 +:temp_w];
assign v307ibus[data_w*2 +:data_w] = c1010obus[data_w*1 +:data_w];
assign c1010ibus[temp_w*2 +:temp_w] = v857obus[temp_w*2 +:temp_w];
assign v857ibus[data_w*2 +:data_w] = c1010obus[data_w*2 +:data_w];
assign c1010ibus[temp_w*3 +:temp_w] = v867obus[temp_w*5 +:temp_w];
assign v867ibus[data_w*5 +:data_w] = c1010obus[data_w*3 +:data_w];
assign c1010ibus[temp_w*4 +:temp_w] = v2162obus[temp_w*1 +:temp_w];
assign v2162ibus[data_w*1 +:data_w] = c1010obus[data_w*4 +:data_w];
assign c1010ibus[temp_w*5 +:temp_w] = v2258obus[temp_w*0 +:temp_w];
assign v2258ibus[data_w*0 +:data_w] = c1010obus[data_w*5 +:data_w];
assign c1011ibus[temp_w*0 +:temp_w] = v250obus[temp_w*5 +:temp_w];
assign v250ibus[data_w*5 +:data_w] = c1011obus[data_w*0 +:data_w];
assign c1011ibus[temp_w*1 +:temp_w] = v308obus[temp_w*2 +:temp_w];
assign v308ibus[data_w*2 +:data_w] = c1011obus[data_w*1 +:data_w];
assign c1011ibus[temp_w*2 +:temp_w] = v858obus[temp_w*2 +:temp_w];
assign v858ibus[data_w*2 +:data_w] = c1011obus[data_w*2 +:data_w];
assign c1011ibus[temp_w*3 +:temp_w] = v868obus[temp_w*5 +:temp_w];
assign v868ibus[data_w*5 +:data_w] = c1011obus[data_w*3 +:data_w];
assign c1011ibus[temp_w*4 +:temp_w] = v2163obus[temp_w*1 +:temp_w];
assign v2163ibus[data_w*1 +:data_w] = c1011obus[data_w*4 +:data_w];
assign c1011ibus[temp_w*5 +:temp_w] = v2259obus[temp_w*0 +:temp_w];
assign v2259ibus[data_w*0 +:data_w] = c1011obus[data_w*5 +:data_w];
assign c1012ibus[temp_w*0 +:temp_w] = v251obus[temp_w*5 +:temp_w];
assign v251ibus[data_w*5 +:data_w] = c1012obus[data_w*0 +:data_w];
assign c1012ibus[temp_w*1 +:temp_w] = v309obus[temp_w*2 +:temp_w];
assign v309ibus[data_w*2 +:data_w] = c1012obus[data_w*1 +:data_w];
assign c1012ibus[temp_w*2 +:temp_w] = v859obus[temp_w*2 +:temp_w];
assign v859ibus[data_w*2 +:data_w] = c1012obus[data_w*2 +:data_w];
assign c1012ibus[temp_w*3 +:temp_w] = v869obus[temp_w*5 +:temp_w];
assign v869ibus[data_w*5 +:data_w] = c1012obus[data_w*3 +:data_w];
assign c1012ibus[temp_w*4 +:temp_w] = v2164obus[temp_w*1 +:temp_w];
assign v2164ibus[data_w*1 +:data_w] = c1012obus[data_w*4 +:data_w];
assign c1012ibus[temp_w*5 +:temp_w] = v2260obus[temp_w*0 +:temp_w];
assign v2260ibus[data_w*0 +:data_w] = c1012obus[data_w*5 +:data_w];
assign c1013ibus[temp_w*0 +:temp_w] = v252obus[temp_w*5 +:temp_w];
assign v252ibus[data_w*5 +:data_w] = c1013obus[data_w*0 +:data_w];
assign c1013ibus[temp_w*1 +:temp_w] = v310obus[temp_w*2 +:temp_w];
assign v310ibus[data_w*2 +:data_w] = c1013obus[data_w*1 +:data_w];
assign c1013ibus[temp_w*2 +:temp_w] = v860obus[temp_w*2 +:temp_w];
assign v860ibus[data_w*2 +:data_w] = c1013obus[data_w*2 +:data_w];
assign c1013ibus[temp_w*3 +:temp_w] = v870obus[temp_w*5 +:temp_w];
assign v870ibus[data_w*5 +:data_w] = c1013obus[data_w*3 +:data_w];
assign c1013ibus[temp_w*4 +:temp_w] = v2165obus[temp_w*1 +:temp_w];
assign v2165ibus[data_w*1 +:data_w] = c1013obus[data_w*4 +:data_w];
assign c1013ibus[temp_w*5 +:temp_w] = v2261obus[temp_w*0 +:temp_w];
assign v2261ibus[data_w*0 +:data_w] = c1013obus[data_w*5 +:data_w];
assign c1014ibus[temp_w*0 +:temp_w] = v253obus[temp_w*5 +:temp_w];
assign v253ibus[data_w*5 +:data_w] = c1014obus[data_w*0 +:data_w];
assign c1014ibus[temp_w*1 +:temp_w] = v311obus[temp_w*2 +:temp_w];
assign v311ibus[data_w*2 +:data_w] = c1014obus[data_w*1 +:data_w];
assign c1014ibus[temp_w*2 +:temp_w] = v861obus[temp_w*2 +:temp_w];
assign v861ibus[data_w*2 +:data_w] = c1014obus[data_w*2 +:data_w];
assign c1014ibus[temp_w*3 +:temp_w] = v871obus[temp_w*5 +:temp_w];
assign v871ibus[data_w*5 +:data_w] = c1014obus[data_w*3 +:data_w];
assign c1014ibus[temp_w*4 +:temp_w] = v2166obus[temp_w*1 +:temp_w];
assign v2166ibus[data_w*1 +:data_w] = c1014obus[data_w*4 +:data_w];
assign c1014ibus[temp_w*5 +:temp_w] = v2262obus[temp_w*0 +:temp_w];
assign v2262ibus[data_w*0 +:data_w] = c1014obus[data_w*5 +:data_w];
assign c1015ibus[temp_w*0 +:temp_w] = v254obus[temp_w*5 +:temp_w];
assign v254ibus[data_w*5 +:data_w] = c1015obus[data_w*0 +:data_w];
assign c1015ibus[temp_w*1 +:temp_w] = v312obus[temp_w*2 +:temp_w];
assign v312ibus[data_w*2 +:data_w] = c1015obus[data_w*1 +:data_w];
assign c1015ibus[temp_w*2 +:temp_w] = v862obus[temp_w*2 +:temp_w];
assign v862ibus[data_w*2 +:data_w] = c1015obus[data_w*2 +:data_w];
assign c1015ibus[temp_w*3 +:temp_w] = v872obus[temp_w*5 +:temp_w];
assign v872ibus[data_w*5 +:data_w] = c1015obus[data_w*3 +:data_w];
assign c1015ibus[temp_w*4 +:temp_w] = v2167obus[temp_w*1 +:temp_w];
assign v2167ibus[data_w*1 +:data_w] = c1015obus[data_w*4 +:data_w];
assign c1015ibus[temp_w*5 +:temp_w] = v2263obus[temp_w*0 +:temp_w];
assign v2263ibus[data_w*0 +:data_w] = c1015obus[data_w*5 +:data_w];
assign c1016ibus[temp_w*0 +:temp_w] = v255obus[temp_w*5 +:temp_w];
assign v255ibus[data_w*5 +:data_w] = c1016obus[data_w*0 +:data_w];
assign c1016ibus[temp_w*1 +:temp_w] = v313obus[temp_w*2 +:temp_w];
assign v313ibus[data_w*2 +:data_w] = c1016obus[data_w*1 +:data_w];
assign c1016ibus[temp_w*2 +:temp_w] = v863obus[temp_w*2 +:temp_w];
assign v863ibus[data_w*2 +:data_w] = c1016obus[data_w*2 +:data_w];
assign c1016ibus[temp_w*3 +:temp_w] = v873obus[temp_w*5 +:temp_w];
assign v873ibus[data_w*5 +:data_w] = c1016obus[data_w*3 +:data_w];
assign c1016ibus[temp_w*4 +:temp_w] = v2168obus[temp_w*1 +:temp_w];
assign v2168ibus[data_w*1 +:data_w] = c1016obus[data_w*4 +:data_w];
assign c1016ibus[temp_w*5 +:temp_w] = v2264obus[temp_w*0 +:temp_w];
assign v2264ibus[data_w*0 +:data_w] = c1016obus[data_w*5 +:data_w];
assign c1017ibus[temp_w*0 +:temp_w] = v256obus[temp_w*5 +:temp_w];
assign v256ibus[data_w*5 +:data_w] = c1017obus[data_w*0 +:data_w];
assign c1017ibus[temp_w*1 +:temp_w] = v314obus[temp_w*2 +:temp_w];
assign v314ibus[data_w*2 +:data_w] = c1017obus[data_w*1 +:data_w];
assign c1017ibus[temp_w*2 +:temp_w] = v768obus[temp_w*2 +:temp_w];
assign v768ibus[data_w*2 +:data_w] = c1017obus[data_w*2 +:data_w];
assign c1017ibus[temp_w*3 +:temp_w] = v874obus[temp_w*5 +:temp_w];
assign v874ibus[data_w*5 +:data_w] = c1017obus[data_w*3 +:data_w];
assign c1017ibus[temp_w*4 +:temp_w] = v2169obus[temp_w*1 +:temp_w];
assign v2169ibus[data_w*1 +:data_w] = c1017obus[data_w*4 +:data_w];
assign c1017ibus[temp_w*5 +:temp_w] = v2265obus[temp_w*0 +:temp_w];
assign v2265ibus[data_w*0 +:data_w] = c1017obus[data_w*5 +:data_w];
assign c1018ibus[temp_w*0 +:temp_w] = v257obus[temp_w*5 +:temp_w];
assign v257ibus[data_w*5 +:data_w] = c1018obus[data_w*0 +:data_w];
assign c1018ibus[temp_w*1 +:temp_w] = v315obus[temp_w*2 +:temp_w];
assign v315ibus[data_w*2 +:data_w] = c1018obus[data_w*1 +:data_w];
assign c1018ibus[temp_w*2 +:temp_w] = v769obus[temp_w*2 +:temp_w];
assign v769ibus[data_w*2 +:data_w] = c1018obus[data_w*2 +:data_w];
assign c1018ibus[temp_w*3 +:temp_w] = v875obus[temp_w*5 +:temp_w];
assign v875ibus[data_w*5 +:data_w] = c1018obus[data_w*3 +:data_w];
assign c1018ibus[temp_w*4 +:temp_w] = v2170obus[temp_w*1 +:temp_w];
assign v2170ibus[data_w*1 +:data_w] = c1018obus[data_w*4 +:data_w];
assign c1018ibus[temp_w*5 +:temp_w] = v2266obus[temp_w*0 +:temp_w];
assign v2266ibus[data_w*0 +:data_w] = c1018obus[data_w*5 +:data_w];
assign c1019ibus[temp_w*0 +:temp_w] = v258obus[temp_w*5 +:temp_w];
assign v258ibus[data_w*5 +:data_w] = c1019obus[data_w*0 +:data_w];
assign c1019ibus[temp_w*1 +:temp_w] = v316obus[temp_w*2 +:temp_w];
assign v316ibus[data_w*2 +:data_w] = c1019obus[data_w*1 +:data_w];
assign c1019ibus[temp_w*2 +:temp_w] = v770obus[temp_w*2 +:temp_w];
assign v770ibus[data_w*2 +:data_w] = c1019obus[data_w*2 +:data_w];
assign c1019ibus[temp_w*3 +:temp_w] = v876obus[temp_w*5 +:temp_w];
assign v876ibus[data_w*5 +:data_w] = c1019obus[data_w*3 +:data_w];
assign c1019ibus[temp_w*4 +:temp_w] = v2171obus[temp_w*1 +:temp_w];
assign v2171ibus[data_w*1 +:data_w] = c1019obus[data_w*4 +:data_w];
assign c1019ibus[temp_w*5 +:temp_w] = v2267obus[temp_w*0 +:temp_w];
assign v2267ibus[data_w*0 +:data_w] = c1019obus[data_w*5 +:data_w];
assign c1020ibus[temp_w*0 +:temp_w] = v259obus[temp_w*5 +:temp_w];
assign v259ibus[data_w*5 +:data_w] = c1020obus[data_w*0 +:data_w];
assign c1020ibus[temp_w*1 +:temp_w] = v317obus[temp_w*2 +:temp_w];
assign v317ibus[data_w*2 +:data_w] = c1020obus[data_w*1 +:data_w];
assign c1020ibus[temp_w*2 +:temp_w] = v771obus[temp_w*2 +:temp_w];
assign v771ibus[data_w*2 +:data_w] = c1020obus[data_w*2 +:data_w];
assign c1020ibus[temp_w*3 +:temp_w] = v877obus[temp_w*5 +:temp_w];
assign v877ibus[data_w*5 +:data_w] = c1020obus[data_w*3 +:data_w];
assign c1020ibus[temp_w*4 +:temp_w] = v2172obus[temp_w*1 +:temp_w];
assign v2172ibus[data_w*1 +:data_w] = c1020obus[data_w*4 +:data_w];
assign c1020ibus[temp_w*5 +:temp_w] = v2268obus[temp_w*0 +:temp_w];
assign v2268ibus[data_w*0 +:data_w] = c1020obus[data_w*5 +:data_w];
assign c1021ibus[temp_w*0 +:temp_w] = v260obus[temp_w*5 +:temp_w];
assign v260ibus[data_w*5 +:data_w] = c1021obus[data_w*0 +:data_w];
assign c1021ibus[temp_w*1 +:temp_w] = v318obus[temp_w*2 +:temp_w];
assign v318ibus[data_w*2 +:data_w] = c1021obus[data_w*1 +:data_w];
assign c1021ibus[temp_w*2 +:temp_w] = v772obus[temp_w*2 +:temp_w];
assign v772ibus[data_w*2 +:data_w] = c1021obus[data_w*2 +:data_w];
assign c1021ibus[temp_w*3 +:temp_w] = v878obus[temp_w*5 +:temp_w];
assign v878ibus[data_w*5 +:data_w] = c1021obus[data_w*3 +:data_w];
assign c1021ibus[temp_w*4 +:temp_w] = v2173obus[temp_w*1 +:temp_w];
assign v2173ibus[data_w*1 +:data_w] = c1021obus[data_w*4 +:data_w];
assign c1021ibus[temp_w*5 +:temp_w] = v2269obus[temp_w*0 +:temp_w];
assign v2269ibus[data_w*0 +:data_w] = c1021obus[data_w*5 +:data_w];
assign c1022ibus[temp_w*0 +:temp_w] = v261obus[temp_w*5 +:temp_w];
assign v261ibus[data_w*5 +:data_w] = c1022obus[data_w*0 +:data_w];
assign c1022ibus[temp_w*1 +:temp_w] = v319obus[temp_w*2 +:temp_w];
assign v319ibus[data_w*2 +:data_w] = c1022obus[data_w*1 +:data_w];
assign c1022ibus[temp_w*2 +:temp_w] = v773obus[temp_w*2 +:temp_w];
assign v773ibus[data_w*2 +:data_w] = c1022obus[data_w*2 +:data_w];
assign c1022ibus[temp_w*3 +:temp_w] = v879obus[temp_w*5 +:temp_w];
assign v879ibus[data_w*5 +:data_w] = c1022obus[data_w*3 +:data_w];
assign c1022ibus[temp_w*4 +:temp_w] = v2174obus[temp_w*1 +:temp_w];
assign v2174ibus[data_w*1 +:data_w] = c1022obus[data_w*4 +:data_w];
assign c1022ibus[temp_w*5 +:temp_w] = v2270obus[temp_w*0 +:temp_w];
assign v2270ibus[data_w*0 +:data_w] = c1022obus[data_w*5 +:data_w];
assign c1023ibus[temp_w*0 +:temp_w] = v262obus[temp_w*5 +:temp_w];
assign v262ibus[data_w*5 +:data_w] = c1023obus[data_w*0 +:data_w];
assign c1023ibus[temp_w*1 +:temp_w] = v320obus[temp_w*2 +:temp_w];
assign v320ibus[data_w*2 +:data_w] = c1023obus[data_w*1 +:data_w];
assign c1023ibus[temp_w*2 +:temp_w] = v774obus[temp_w*2 +:temp_w];
assign v774ibus[data_w*2 +:data_w] = c1023obus[data_w*2 +:data_w];
assign c1023ibus[temp_w*3 +:temp_w] = v880obus[temp_w*5 +:temp_w];
assign v880ibus[data_w*5 +:data_w] = c1023obus[data_w*3 +:data_w];
assign c1023ibus[temp_w*4 +:temp_w] = v2175obus[temp_w*1 +:temp_w];
assign v2175ibus[data_w*1 +:data_w] = c1023obus[data_w*4 +:data_w];
assign c1023ibus[temp_w*5 +:temp_w] = v2271obus[temp_w*0 +:temp_w];
assign v2271ibus[data_w*0 +:data_w] = c1023obus[data_w*5 +:data_w];
assign c1024ibus[temp_w*0 +:temp_w] = v263obus[temp_w*5 +:temp_w];
assign v263ibus[data_w*5 +:data_w] = c1024obus[data_w*0 +:data_w];
assign c1024ibus[temp_w*1 +:temp_w] = v321obus[temp_w*2 +:temp_w];
assign v321ibus[data_w*2 +:data_w] = c1024obus[data_w*1 +:data_w];
assign c1024ibus[temp_w*2 +:temp_w] = v775obus[temp_w*2 +:temp_w];
assign v775ibus[data_w*2 +:data_w] = c1024obus[data_w*2 +:data_w];
assign c1024ibus[temp_w*3 +:temp_w] = v881obus[temp_w*5 +:temp_w];
assign v881ibus[data_w*5 +:data_w] = c1024obus[data_w*3 +:data_w];
assign c1024ibus[temp_w*4 +:temp_w] = v2176obus[temp_w*1 +:temp_w];
assign v2176ibus[data_w*1 +:data_w] = c1024obus[data_w*4 +:data_w];
assign c1024ibus[temp_w*5 +:temp_w] = v2272obus[temp_w*0 +:temp_w];
assign v2272ibus[data_w*0 +:data_w] = c1024obus[data_w*5 +:data_w];
assign c1025ibus[temp_w*0 +:temp_w] = v264obus[temp_w*5 +:temp_w];
assign v264ibus[data_w*5 +:data_w] = c1025obus[data_w*0 +:data_w];
assign c1025ibus[temp_w*1 +:temp_w] = v322obus[temp_w*2 +:temp_w];
assign v322ibus[data_w*2 +:data_w] = c1025obus[data_w*1 +:data_w];
assign c1025ibus[temp_w*2 +:temp_w] = v776obus[temp_w*2 +:temp_w];
assign v776ibus[data_w*2 +:data_w] = c1025obus[data_w*2 +:data_w];
assign c1025ibus[temp_w*3 +:temp_w] = v882obus[temp_w*5 +:temp_w];
assign v882ibus[data_w*5 +:data_w] = c1025obus[data_w*3 +:data_w];
assign c1025ibus[temp_w*4 +:temp_w] = v2177obus[temp_w*1 +:temp_w];
assign v2177ibus[data_w*1 +:data_w] = c1025obus[data_w*4 +:data_w];
assign c1025ibus[temp_w*5 +:temp_w] = v2273obus[temp_w*0 +:temp_w];
assign v2273ibus[data_w*0 +:data_w] = c1025obus[data_w*5 +:data_w];
assign c1026ibus[temp_w*0 +:temp_w] = v265obus[temp_w*5 +:temp_w];
assign v265ibus[data_w*5 +:data_w] = c1026obus[data_w*0 +:data_w];
assign c1026ibus[temp_w*1 +:temp_w] = v323obus[temp_w*2 +:temp_w];
assign v323ibus[data_w*2 +:data_w] = c1026obus[data_w*1 +:data_w];
assign c1026ibus[temp_w*2 +:temp_w] = v777obus[temp_w*2 +:temp_w];
assign v777ibus[data_w*2 +:data_w] = c1026obus[data_w*2 +:data_w];
assign c1026ibus[temp_w*3 +:temp_w] = v883obus[temp_w*5 +:temp_w];
assign v883ibus[data_w*5 +:data_w] = c1026obus[data_w*3 +:data_w];
assign c1026ibus[temp_w*4 +:temp_w] = v2178obus[temp_w*1 +:temp_w];
assign v2178ibus[data_w*1 +:data_w] = c1026obus[data_w*4 +:data_w];
assign c1026ibus[temp_w*5 +:temp_w] = v2274obus[temp_w*0 +:temp_w];
assign v2274ibus[data_w*0 +:data_w] = c1026obus[data_w*5 +:data_w];
assign c1027ibus[temp_w*0 +:temp_w] = v266obus[temp_w*5 +:temp_w];
assign v266ibus[data_w*5 +:data_w] = c1027obus[data_w*0 +:data_w];
assign c1027ibus[temp_w*1 +:temp_w] = v324obus[temp_w*2 +:temp_w];
assign v324ibus[data_w*2 +:data_w] = c1027obus[data_w*1 +:data_w];
assign c1027ibus[temp_w*2 +:temp_w] = v778obus[temp_w*2 +:temp_w];
assign v778ibus[data_w*2 +:data_w] = c1027obus[data_w*2 +:data_w];
assign c1027ibus[temp_w*3 +:temp_w] = v884obus[temp_w*5 +:temp_w];
assign v884ibus[data_w*5 +:data_w] = c1027obus[data_w*3 +:data_w];
assign c1027ibus[temp_w*4 +:temp_w] = v2179obus[temp_w*1 +:temp_w];
assign v2179ibus[data_w*1 +:data_w] = c1027obus[data_w*4 +:data_w];
assign c1027ibus[temp_w*5 +:temp_w] = v2275obus[temp_w*0 +:temp_w];
assign v2275ibus[data_w*0 +:data_w] = c1027obus[data_w*5 +:data_w];
assign c1028ibus[temp_w*0 +:temp_w] = v267obus[temp_w*5 +:temp_w];
assign v267ibus[data_w*5 +:data_w] = c1028obus[data_w*0 +:data_w];
assign c1028ibus[temp_w*1 +:temp_w] = v325obus[temp_w*2 +:temp_w];
assign v325ibus[data_w*2 +:data_w] = c1028obus[data_w*1 +:data_w];
assign c1028ibus[temp_w*2 +:temp_w] = v779obus[temp_w*2 +:temp_w];
assign v779ibus[data_w*2 +:data_w] = c1028obus[data_w*2 +:data_w];
assign c1028ibus[temp_w*3 +:temp_w] = v885obus[temp_w*5 +:temp_w];
assign v885ibus[data_w*5 +:data_w] = c1028obus[data_w*3 +:data_w];
assign c1028ibus[temp_w*4 +:temp_w] = v2180obus[temp_w*1 +:temp_w];
assign v2180ibus[data_w*1 +:data_w] = c1028obus[data_w*4 +:data_w];
assign c1028ibus[temp_w*5 +:temp_w] = v2276obus[temp_w*0 +:temp_w];
assign v2276ibus[data_w*0 +:data_w] = c1028obus[data_w*5 +:data_w];
assign c1029ibus[temp_w*0 +:temp_w] = v268obus[temp_w*5 +:temp_w];
assign v268ibus[data_w*5 +:data_w] = c1029obus[data_w*0 +:data_w];
assign c1029ibus[temp_w*1 +:temp_w] = v326obus[temp_w*2 +:temp_w];
assign v326ibus[data_w*2 +:data_w] = c1029obus[data_w*1 +:data_w];
assign c1029ibus[temp_w*2 +:temp_w] = v780obus[temp_w*2 +:temp_w];
assign v780ibus[data_w*2 +:data_w] = c1029obus[data_w*2 +:data_w];
assign c1029ibus[temp_w*3 +:temp_w] = v886obus[temp_w*5 +:temp_w];
assign v886ibus[data_w*5 +:data_w] = c1029obus[data_w*3 +:data_w];
assign c1029ibus[temp_w*4 +:temp_w] = v2181obus[temp_w*1 +:temp_w];
assign v2181ibus[data_w*1 +:data_w] = c1029obus[data_w*4 +:data_w];
assign c1029ibus[temp_w*5 +:temp_w] = v2277obus[temp_w*0 +:temp_w];
assign v2277ibus[data_w*0 +:data_w] = c1029obus[data_w*5 +:data_w];
assign c1030ibus[temp_w*0 +:temp_w] = v269obus[temp_w*5 +:temp_w];
assign v269ibus[data_w*5 +:data_w] = c1030obus[data_w*0 +:data_w];
assign c1030ibus[temp_w*1 +:temp_w] = v327obus[temp_w*2 +:temp_w];
assign v327ibus[data_w*2 +:data_w] = c1030obus[data_w*1 +:data_w];
assign c1030ibus[temp_w*2 +:temp_w] = v781obus[temp_w*2 +:temp_w];
assign v781ibus[data_w*2 +:data_w] = c1030obus[data_w*2 +:data_w];
assign c1030ibus[temp_w*3 +:temp_w] = v887obus[temp_w*5 +:temp_w];
assign v887ibus[data_w*5 +:data_w] = c1030obus[data_w*3 +:data_w];
assign c1030ibus[temp_w*4 +:temp_w] = v2182obus[temp_w*1 +:temp_w];
assign v2182ibus[data_w*1 +:data_w] = c1030obus[data_w*4 +:data_w];
assign c1030ibus[temp_w*5 +:temp_w] = v2278obus[temp_w*0 +:temp_w];
assign v2278ibus[data_w*0 +:data_w] = c1030obus[data_w*5 +:data_w];
assign c1031ibus[temp_w*0 +:temp_w] = v270obus[temp_w*5 +:temp_w];
assign v270ibus[data_w*5 +:data_w] = c1031obus[data_w*0 +:data_w];
assign c1031ibus[temp_w*1 +:temp_w] = v328obus[temp_w*2 +:temp_w];
assign v328ibus[data_w*2 +:data_w] = c1031obus[data_w*1 +:data_w];
assign c1031ibus[temp_w*2 +:temp_w] = v782obus[temp_w*2 +:temp_w];
assign v782ibus[data_w*2 +:data_w] = c1031obus[data_w*2 +:data_w];
assign c1031ibus[temp_w*3 +:temp_w] = v888obus[temp_w*5 +:temp_w];
assign v888ibus[data_w*5 +:data_w] = c1031obus[data_w*3 +:data_w];
assign c1031ibus[temp_w*4 +:temp_w] = v2183obus[temp_w*1 +:temp_w];
assign v2183ibus[data_w*1 +:data_w] = c1031obus[data_w*4 +:data_w];
assign c1031ibus[temp_w*5 +:temp_w] = v2279obus[temp_w*0 +:temp_w];
assign v2279ibus[data_w*0 +:data_w] = c1031obus[data_w*5 +:data_w];
assign c1032ibus[temp_w*0 +:temp_w] = v271obus[temp_w*5 +:temp_w];
assign v271ibus[data_w*5 +:data_w] = c1032obus[data_w*0 +:data_w];
assign c1032ibus[temp_w*1 +:temp_w] = v329obus[temp_w*2 +:temp_w];
assign v329ibus[data_w*2 +:data_w] = c1032obus[data_w*1 +:data_w];
assign c1032ibus[temp_w*2 +:temp_w] = v783obus[temp_w*2 +:temp_w];
assign v783ibus[data_w*2 +:data_w] = c1032obus[data_w*2 +:data_w];
assign c1032ibus[temp_w*3 +:temp_w] = v889obus[temp_w*5 +:temp_w];
assign v889ibus[data_w*5 +:data_w] = c1032obus[data_w*3 +:data_w];
assign c1032ibus[temp_w*4 +:temp_w] = v2184obus[temp_w*1 +:temp_w];
assign v2184ibus[data_w*1 +:data_w] = c1032obus[data_w*4 +:data_w];
assign c1032ibus[temp_w*5 +:temp_w] = v2280obus[temp_w*0 +:temp_w];
assign v2280ibus[data_w*0 +:data_w] = c1032obus[data_w*5 +:data_w];
assign c1033ibus[temp_w*0 +:temp_w] = v272obus[temp_w*5 +:temp_w];
assign v272ibus[data_w*5 +:data_w] = c1033obus[data_w*0 +:data_w];
assign c1033ibus[temp_w*1 +:temp_w] = v330obus[temp_w*2 +:temp_w];
assign v330ibus[data_w*2 +:data_w] = c1033obus[data_w*1 +:data_w];
assign c1033ibus[temp_w*2 +:temp_w] = v784obus[temp_w*2 +:temp_w];
assign v784ibus[data_w*2 +:data_w] = c1033obus[data_w*2 +:data_w];
assign c1033ibus[temp_w*3 +:temp_w] = v890obus[temp_w*5 +:temp_w];
assign v890ibus[data_w*5 +:data_w] = c1033obus[data_w*3 +:data_w];
assign c1033ibus[temp_w*4 +:temp_w] = v2185obus[temp_w*1 +:temp_w];
assign v2185ibus[data_w*1 +:data_w] = c1033obus[data_w*4 +:data_w];
assign c1033ibus[temp_w*5 +:temp_w] = v2281obus[temp_w*0 +:temp_w];
assign v2281ibus[data_w*0 +:data_w] = c1033obus[data_w*5 +:data_w];
assign c1034ibus[temp_w*0 +:temp_w] = v273obus[temp_w*5 +:temp_w];
assign v273ibus[data_w*5 +:data_w] = c1034obus[data_w*0 +:data_w];
assign c1034ibus[temp_w*1 +:temp_w] = v331obus[temp_w*2 +:temp_w];
assign v331ibus[data_w*2 +:data_w] = c1034obus[data_w*1 +:data_w];
assign c1034ibus[temp_w*2 +:temp_w] = v785obus[temp_w*2 +:temp_w];
assign v785ibus[data_w*2 +:data_w] = c1034obus[data_w*2 +:data_w];
assign c1034ibus[temp_w*3 +:temp_w] = v891obus[temp_w*5 +:temp_w];
assign v891ibus[data_w*5 +:data_w] = c1034obus[data_w*3 +:data_w];
assign c1034ibus[temp_w*4 +:temp_w] = v2186obus[temp_w*1 +:temp_w];
assign v2186ibus[data_w*1 +:data_w] = c1034obus[data_w*4 +:data_w];
assign c1034ibus[temp_w*5 +:temp_w] = v2282obus[temp_w*0 +:temp_w];
assign v2282ibus[data_w*0 +:data_w] = c1034obus[data_w*5 +:data_w];
assign c1035ibus[temp_w*0 +:temp_w] = v274obus[temp_w*5 +:temp_w];
assign v274ibus[data_w*5 +:data_w] = c1035obus[data_w*0 +:data_w];
assign c1035ibus[temp_w*1 +:temp_w] = v332obus[temp_w*2 +:temp_w];
assign v332ibus[data_w*2 +:data_w] = c1035obus[data_w*1 +:data_w];
assign c1035ibus[temp_w*2 +:temp_w] = v786obus[temp_w*2 +:temp_w];
assign v786ibus[data_w*2 +:data_w] = c1035obus[data_w*2 +:data_w];
assign c1035ibus[temp_w*3 +:temp_w] = v892obus[temp_w*5 +:temp_w];
assign v892ibus[data_w*5 +:data_w] = c1035obus[data_w*3 +:data_w];
assign c1035ibus[temp_w*4 +:temp_w] = v2187obus[temp_w*1 +:temp_w];
assign v2187ibus[data_w*1 +:data_w] = c1035obus[data_w*4 +:data_w];
assign c1035ibus[temp_w*5 +:temp_w] = v2283obus[temp_w*0 +:temp_w];
assign v2283ibus[data_w*0 +:data_w] = c1035obus[data_w*5 +:data_w];
assign c1036ibus[temp_w*0 +:temp_w] = v275obus[temp_w*5 +:temp_w];
assign v275ibus[data_w*5 +:data_w] = c1036obus[data_w*0 +:data_w];
assign c1036ibus[temp_w*1 +:temp_w] = v333obus[temp_w*2 +:temp_w];
assign v333ibus[data_w*2 +:data_w] = c1036obus[data_w*1 +:data_w];
assign c1036ibus[temp_w*2 +:temp_w] = v787obus[temp_w*2 +:temp_w];
assign v787ibus[data_w*2 +:data_w] = c1036obus[data_w*2 +:data_w];
assign c1036ibus[temp_w*3 +:temp_w] = v893obus[temp_w*5 +:temp_w];
assign v893ibus[data_w*5 +:data_w] = c1036obus[data_w*3 +:data_w];
assign c1036ibus[temp_w*4 +:temp_w] = v2188obus[temp_w*1 +:temp_w];
assign v2188ibus[data_w*1 +:data_w] = c1036obus[data_w*4 +:data_w];
assign c1036ibus[temp_w*5 +:temp_w] = v2284obus[temp_w*0 +:temp_w];
assign v2284ibus[data_w*0 +:data_w] = c1036obus[data_w*5 +:data_w];
assign c1037ibus[temp_w*0 +:temp_w] = v276obus[temp_w*5 +:temp_w];
assign v276ibus[data_w*5 +:data_w] = c1037obus[data_w*0 +:data_w];
assign c1037ibus[temp_w*1 +:temp_w] = v334obus[temp_w*2 +:temp_w];
assign v334ibus[data_w*2 +:data_w] = c1037obus[data_w*1 +:data_w];
assign c1037ibus[temp_w*2 +:temp_w] = v788obus[temp_w*2 +:temp_w];
assign v788ibus[data_w*2 +:data_w] = c1037obus[data_w*2 +:data_w];
assign c1037ibus[temp_w*3 +:temp_w] = v894obus[temp_w*5 +:temp_w];
assign v894ibus[data_w*5 +:data_w] = c1037obus[data_w*3 +:data_w];
assign c1037ibus[temp_w*4 +:temp_w] = v2189obus[temp_w*1 +:temp_w];
assign v2189ibus[data_w*1 +:data_w] = c1037obus[data_w*4 +:data_w];
assign c1037ibus[temp_w*5 +:temp_w] = v2285obus[temp_w*0 +:temp_w];
assign v2285ibus[data_w*0 +:data_w] = c1037obus[data_w*5 +:data_w];
assign c1038ibus[temp_w*0 +:temp_w] = v277obus[temp_w*5 +:temp_w];
assign v277ibus[data_w*5 +:data_w] = c1038obus[data_w*0 +:data_w];
assign c1038ibus[temp_w*1 +:temp_w] = v335obus[temp_w*2 +:temp_w];
assign v335ibus[data_w*2 +:data_w] = c1038obus[data_w*1 +:data_w];
assign c1038ibus[temp_w*2 +:temp_w] = v789obus[temp_w*2 +:temp_w];
assign v789ibus[data_w*2 +:data_w] = c1038obus[data_w*2 +:data_w];
assign c1038ibus[temp_w*3 +:temp_w] = v895obus[temp_w*5 +:temp_w];
assign v895ibus[data_w*5 +:data_w] = c1038obus[data_w*3 +:data_w];
assign c1038ibus[temp_w*4 +:temp_w] = v2190obus[temp_w*1 +:temp_w];
assign v2190ibus[data_w*1 +:data_w] = c1038obus[data_w*4 +:data_w];
assign c1038ibus[temp_w*5 +:temp_w] = v2286obus[temp_w*0 +:temp_w];
assign v2286ibus[data_w*0 +:data_w] = c1038obus[data_w*5 +:data_w];
assign c1039ibus[temp_w*0 +:temp_w] = v278obus[temp_w*5 +:temp_w];
assign v278ibus[data_w*5 +:data_w] = c1039obus[data_w*0 +:data_w];
assign c1039ibus[temp_w*1 +:temp_w] = v336obus[temp_w*2 +:temp_w];
assign v336ibus[data_w*2 +:data_w] = c1039obus[data_w*1 +:data_w];
assign c1039ibus[temp_w*2 +:temp_w] = v790obus[temp_w*2 +:temp_w];
assign v790ibus[data_w*2 +:data_w] = c1039obus[data_w*2 +:data_w];
assign c1039ibus[temp_w*3 +:temp_w] = v896obus[temp_w*5 +:temp_w];
assign v896ibus[data_w*5 +:data_w] = c1039obus[data_w*3 +:data_w];
assign c1039ibus[temp_w*4 +:temp_w] = v2191obus[temp_w*1 +:temp_w];
assign v2191ibus[data_w*1 +:data_w] = c1039obus[data_w*4 +:data_w];
assign c1039ibus[temp_w*5 +:temp_w] = v2287obus[temp_w*0 +:temp_w];
assign v2287ibus[data_w*0 +:data_w] = c1039obus[data_w*5 +:data_w];
assign c1040ibus[temp_w*0 +:temp_w] = v279obus[temp_w*5 +:temp_w];
assign v279ibus[data_w*5 +:data_w] = c1040obus[data_w*0 +:data_w];
assign c1040ibus[temp_w*1 +:temp_w] = v337obus[temp_w*2 +:temp_w];
assign v337ibus[data_w*2 +:data_w] = c1040obus[data_w*1 +:data_w];
assign c1040ibus[temp_w*2 +:temp_w] = v791obus[temp_w*2 +:temp_w];
assign v791ibus[data_w*2 +:data_w] = c1040obus[data_w*2 +:data_w];
assign c1040ibus[temp_w*3 +:temp_w] = v897obus[temp_w*5 +:temp_w];
assign v897ibus[data_w*5 +:data_w] = c1040obus[data_w*3 +:data_w];
assign c1040ibus[temp_w*4 +:temp_w] = v2192obus[temp_w*1 +:temp_w];
assign v2192ibus[data_w*1 +:data_w] = c1040obus[data_w*4 +:data_w];
assign c1040ibus[temp_w*5 +:temp_w] = v2288obus[temp_w*0 +:temp_w];
assign v2288ibus[data_w*0 +:data_w] = c1040obus[data_w*5 +:data_w];
assign c1041ibus[temp_w*0 +:temp_w] = v280obus[temp_w*5 +:temp_w];
assign v280ibus[data_w*5 +:data_w] = c1041obus[data_w*0 +:data_w];
assign c1041ibus[temp_w*1 +:temp_w] = v338obus[temp_w*2 +:temp_w];
assign v338ibus[data_w*2 +:data_w] = c1041obus[data_w*1 +:data_w];
assign c1041ibus[temp_w*2 +:temp_w] = v792obus[temp_w*2 +:temp_w];
assign v792ibus[data_w*2 +:data_w] = c1041obus[data_w*2 +:data_w];
assign c1041ibus[temp_w*3 +:temp_w] = v898obus[temp_w*5 +:temp_w];
assign v898ibus[data_w*5 +:data_w] = c1041obus[data_w*3 +:data_w];
assign c1041ibus[temp_w*4 +:temp_w] = v2193obus[temp_w*1 +:temp_w];
assign v2193ibus[data_w*1 +:data_w] = c1041obus[data_w*4 +:data_w];
assign c1041ibus[temp_w*5 +:temp_w] = v2289obus[temp_w*0 +:temp_w];
assign v2289ibus[data_w*0 +:data_w] = c1041obus[data_w*5 +:data_w];
assign c1042ibus[temp_w*0 +:temp_w] = v281obus[temp_w*5 +:temp_w];
assign v281ibus[data_w*5 +:data_w] = c1042obus[data_w*0 +:data_w];
assign c1042ibus[temp_w*1 +:temp_w] = v339obus[temp_w*2 +:temp_w];
assign v339ibus[data_w*2 +:data_w] = c1042obus[data_w*1 +:data_w];
assign c1042ibus[temp_w*2 +:temp_w] = v793obus[temp_w*2 +:temp_w];
assign v793ibus[data_w*2 +:data_w] = c1042obus[data_w*2 +:data_w];
assign c1042ibus[temp_w*3 +:temp_w] = v899obus[temp_w*5 +:temp_w];
assign v899ibus[data_w*5 +:data_w] = c1042obus[data_w*3 +:data_w];
assign c1042ibus[temp_w*4 +:temp_w] = v2194obus[temp_w*1 +:temp_w];
assign v2194ibus[data_w*1 +:data_w] = c1042obus[data_w*4 +:data_w];
assign c1042ibus[temp_w*5 +:temp_w] = v2290obus[temp_w*0 +:temp_w];
assign v2290ibus[data_w*0 +:data_w] = c1042obus[data_w*5 +:data_w];
assign c1043ibus[temp_w*0 +:temp_w] = v282obus[temp_w*5 +:temp_w];
assign v282ibus[data_w*5 +:data_w] = c1043obus[data_w*0 +:data_w];
assign c1043ibus[temp_w*1 +:temp_w] = v340obus[temp_w*2 +:temp_w];
assign v340ibus[data_w*2 +:data_w] = c1043obus[data_w*1 +:data_w];
assign c1043ibus[temp_w*2 +:temp_w] = v794obus[temp_w*2 +:temp_w];
assign v794ibus[data_w*2 +:data_w] = c1043obus[data_w*2 +:data_w];
assign c1043ibus[temp_w*3 +:temp_w] = v900obus[temp_w*5 +:temp_w];
assign v900ibus[data_w*5 +:data_w] = c1043obus[data_w*3 +:data_w];
assign c1043ibus[temp_w*4 +:temp_w] = v2195obus[temp_w*1 +:temp_w];
assign v2195ibus[data_w*1 +:data_w] = c1043obus[data_w*4 +:data_w];
assign c1043ibus[temp_w*5 +:temp_w] = v2291obus[temp_w*0 +:temp_w];
assign v2291ibus[data_w*0 +:data_w] = c1043obus[data_w*5 +:data_w];
assign c1044ibus[temp_w*0 +:temp_w] = v283obus[temp_w*5 +:temp_w];
assign v283ibus[data_w*5 +:data_w] = c1044obus[data_w*0 +:data_w];
assign c1044ibus[temp_w*1 +:temp_w] = v341obus[temp_w*2 +:temp_w];
assign v341ibus[data_w*2 +:data_w] = c1044obus[data_w*1 +:data_w];
assign c1044ibus[temp_w*2 +:temp_w] = v795obus[temp_w*2 +:temp_w];
assign v795ibus[data_w*2 +:data_w] = c1044obus[data_w*2 +:data_w];
assign c1044ibus[temp_w*3 +:temp_w] = v901obus[temp_w*5 +:temp_w];
assign v901ibus[data_w*5 +:data_w] = c1044obus[data_w*3 +:data_w];
assign c1044ibus[temp_w*4 +:temp_w] = v2196obus[temp_w*1 +:temp_w];
assign v2196ibus[data_w*1 +:data_w] = c1044obus[data_w*4 +:data_w];
assign c1044ibus[temp_w*5 +:temp_w] = v2292obus[temp_w*0 +:temp_w];
assign v2292ibus[data_w*0 +:data_w] = c1044obus[data_w*5 +:data_w];
assign c1045ibus[temp_w*0 +:temp_w] = v284obus[temp_w*5 +:temp_w];
assign v284ibus[data_w*5 +:data_w] = c1045obus[data_w*0 +:data_w];
assign c1045ibus[temp_w*1 +:temp_w] = v342obus[temp_w*2 +:temp_w];
assign v342ibus[data_w*2 +:data_w] = c1045obus[data_w*1 +:data_w];
assign c1045ibus[temp_w*2 +:temp_w] = v796obus[temp_w*2 +:temp_w];
assign v796ibus[data_w*2 +:data_w] = c1045obus[data_w*2 +:data_w];
assign c1045ibus[temp_w*3 +:temp_w] = v902obus[temp_w*5 +:temp_w];
assign v902ibus[data_w*5 +:data_w] = c1045obus[data_w*3 +:data_w];
assign c1045ibus[temp_w*4 +:temp_w] = v2197obus[temp_w*1 +:temp_w];
assign v2197ibus[data_w*1 +:data_w] = c1045obus[data_w*4 +:data_w];
assign c1045ibus[temp_w*5 +:temp_w] = v2293obus[temp_w*0 +:temp_w];
assign v2293ibus[data_w*0 +:data_w] = c1045obus[data_w*5 +:data_w];
assign c1046ibus[temp_w*0 +:temp_w] = v285obus[temp_w*5 +:temp_w];
assign v285ibus[data_w*5 +:data_w] = c1046obus[data_w*0 +:data_w];
assign c1046ibus[temp_w*1 +:temp_w] = v343obus[temp_w*2 +:temp_w];
assign v343ibus[data_w*2 +:data_w] = c1046obus[data_w*1 +:data_w];
assign c1046ibus[temp_w*2 +:temp_w] = v797obus[temp_w*2 +:temp_w];
assign v797ibus[data_w*2 +:data_w] = c1046obus[data_w*2 +:data_w];
assign c1046ibus[temp_w*3 +:temp_w] = v903obus[temp_w*5 +:temp_w];
assign v903ibus[data_w*5 +:data_w] = c1046obus[data_w*3 +:data_w];
assign c1046ibus[temp_w*4 +:temp_w] = v2198obus[temp_w*1 +:temp_w];
assign v2198ibus[data_w*1 +:data_w] = c1046obus[data_w*4 +:data_w];
assign c1046ibus[temp_w*5 +:temp_w] = v2294obus[temp_w*0 +:temp_w];
assign v2294ibus[data_w*0 +:data_w] = c1046obus[data_w*5 +:data_w];
assign c1047ibus[temp_w*0 +:temp_w] = v286obus[temp_w*5 +:temp_w];
assign v286ibus[data_w*5 +:data_w] = c1047obus[data_w*0 +:data_w];
assign c1047ibus[temp_w*1 +:temp_w] = v344obus[temp_w*2 +:temp_w];
assign v344ibus[data_w*2 +:data_w] = c1047obus[data_w*1 +:data_w];
assign c1047ibus[temp_w*2 +:temp_w] = v798obus[temp_w*2 +:temp_w];
assign v798ibus[data_w*2 +:data_w] = c1047obus[data_w*2 +:data_w];
assign c1047ibus[temp_w*3 +:temp_w] = v904obus[temp_w*5 +:temp_w];
assign v904ibus[data_w*5 +:data_w] = c1047obus[data_w*3 +:data_w];
assign c1047ibus[temp_w*4 +:temp_w] = v2199obus[temp_w*1 +:temp_w];
assign v2199ibus[data_w*1 +:data_w] = c1047obus[data_w*4 +:data_w];
assign c1047ibus[temp_w*5 +:temp_w] = v2295obus[temp_w*0 +:temp_w];
assign v2295ibus[data_w*0 +:data_w] = c1047obus[data_w*5 +:data_w];
assign c1048ibus[temp_w*0 +:temp_w] = v287obus[temp_w*5 +:temp_w];
assign v287ibus[data_w*5 +:data_w] = c1048obus[data_w*0 +:data_w];
assign c1048ibus[temp_w*1 +:temp_w] = v345obus[temp_w*2 +:temp_w];
assign v345ibus[data_w*2 +:data_w] = c1048obus[data_w*1 +:data_w];
assign c1048ibus[temp_w*2 +:temp_w] = v799obus[temp_w*2 +:temp_w];
assign v799ibus[data_w*2 +:data_w] = c1048obus[data_w*2 +:data_w];
assign c1048ibus[temp_w*3 +:temp_w] = v905obus[temp_w*5 +:temp_w];
assign v905ibus[data_w*5 +:data_w] = c1048obus[data_w*3 +:data_w];
assign c1048ibus[temp_w*4 +:temp_w] = v2200obus[temp_w*1 +:temp_w];
assign v2200ibus[data_w*1 +:data_w] = c1048obus[data_w*4 +:data_w];
assign c1048ibus[temp_w*5 +:temp_w] = v2296obus[temp_w*0 +:temp_w];
assign v2296ibus[data_w*0 +:data_w] = c1048obus[data_w*5 +:data_w];
assign c1049ibus[temp_w*0 +:temp_w] = v192obus[temp_w*5 +:temp_w];
assign v192ibus[data_w*5 +:data_w] = c1049obus[data_w*0 +:data_w];
assign c1049ibus[temp_w*1 +:temp_w] = v346obus[temp_w*2 +:temp_w];
assign v346ibus[data_w*2 +:data_w] = c1049obus[data_w*1 +:data_w];
assign c1049ibus[temp_w*2 +:temp_w] = v800obus[temp_w*2 +:temp_w];
assign v800ibus[data_w*2 +:data_w] = c1049obus[data_w*2 +:data_w];
assign c1049ibus[temp_w*3 +:temp_w] = v906obus[temp_w*5 +:temp_w];
assign v906ibus[data_w*5 +:data_w] = c1049obus[data_w*3 +:data_w];
assign c1049ibus[temp_w*4 +:temp_w] = v2201obus[temp_w*1 +:temp_w];
assign v2201ibus[data_w*1 +:data_w] = c1049obus[data_w*4 +:data_w];
assign c1049ibus[temp_w*5 +:temp_w] = v2297obus[temp_w*0 +:temp_w];
assign v2297ibus[data_w*0 +:data_w] = c1049obus[data_w*5 +:data_w];
assign c1050ibus[temp_w*0 +:temp_w] = v193obus[temp_w*5 +:temp_w];
assign v193ibus[data_w*5 +:data_w] = c1050obus[data_w*0 +:data_w];
assign c1050ibus[temp_w*1 +:temp_w] = v347obus[temp_w*2 +:temp_w];
assign v347ibus[data_w*2 +:data_w] = c1050obus[data_w*1 +:data_w];
assign c1050ibus[temp_w*2 +:temp_w] = v801obus[temp_w*2 +:temp_w];
assign v801ibus[data_w*2 +:data_w] = c1050obus[data_w*2 +:data_w];
assign c1050ibus[temp_w*3 +:temp_w] = v907obus[temp_w*5 +:temp_w];
assign v907ibus[data_w*5 +:data_w] = c1050obus[data_w*3 +:data_w];
assign c1050ibus[temp_w*4 +:temp_w] = v2202obus[temp_w*1 +:temp_w];
assign v2202ibus[data_w*1 +:data_w] = c1050obus[data_w*4 +:data_w];
assign c1050ibus[temp_w*5 +:temp_w] = v2298obus[temp_w*0 +:temp_w];
assign v2298ibus[data_w*0 +:data_w] = c1050obus[data_w*5 +:data_w];
assign c1051ibus[temp_w*0 +:temp_w] = v194obus[temp_w*5 +:temp_w];
assign v194ibus[data_w*5 +:data_w] = c1051obus[data_w*0 +:data_w];
assign c1051ibus[temp_w*1 +:temp_w] = v348obus[temp_w*2 +:temp_w];
assign v348ibus[data_w*2 +:data_w] = c1051obus[data_w*1 +:data_w];
assign c1051ibus[temp_w*2 +:temp_w] = v802obus[temp_w*2 +:temp_w];
assign v802ibus[data_w*2 +:data_w] = c1051obus[data_w*2 +:data_w];
assign c1051ibus[temp_w*3 +:temp_w] = v908obus[temp_w*5 +:temp_w];
assign v908ibus[data_w*5 +:data_w] = c1051obus[data_w*3 +:data_w];
assign c1051ibus[temp_w*4 +:temp_w] = v2203obus[temp_w*1 +:temp_w];
assign v2203ibus[data_w*1 +:data_w] = c1051obus[data_w*4 +:data_w];
assign c1051ibus[temp_w*5 +:temp_w] = v2299obus[temp_w*0 +:temp_w];
assign v2299ibus[data_w*0 +:data_w] = c1051obus[data_w*5 +:data_w];
assign c1052ibus[temp_w*0 +:temp_w] = v195obus[temp_w*5 +:temp_w];
assign v195ibus[data_w*5 +:data_w] = c1052obus[data_w*0 +:data_w];
assign c1052ibus[temp_w*1 +:temp_w] = v349obus[temp_w*2 +:temp_w];
assign v349ibus[data_w*2 +:data_w] = c1052obus[data_w*1 +:data_w];
assign c1052ibus[temp_w*2 +:temp_w] = v803obus[temp_w*2 +:temp_w];
assign v803ibus[data_w*2 +:data_w] = c1052obus[data_w*2 +:data_w];
assign c1052ibus[temp_w*3 +:temp_w] = v909obus[temp_w*5 +:temp_w];
assign v909ibus[data_w*5 +:data_w] = c1052obus[data_w*3 +:data_w];
assign c1052ibus[temp_w*4 +:temp_w] = v2204obus[temp_w*1 +:temp_w];
assign v2204ibus[data_w*1 +:data_w] = c1052obus[data_w*4 +:data_w];
assign c1052ibus[temp_w*5 +:temp_w] = v2300obus[temp_w*0 +:temp_w];
assign v2300ibus[data_w*0 +:data_w] = c1052obus[data_w*5 +:data_w];
assign c1053ibus[temp_w*0 +:temp_w] = v196obus[temp_w*5 +:temp_w];
assign v196ibus[data_w*5 +:data_w] = c1053obus[data_w*0 +:data_w];
assign c1053ibus[temp_w*1 +:temp_w] = v350obus[temp_w*2 +:temp_w];
assign v350ibus[data_w*2 +:data_w] = c1053obus[data_w*1 +:data_w];
assign c1053ibus[temp_w*2 +:temp_w] = v804obus[temp_w*2 +:temp_w];
assign v804ibus[data_w*2 +:data_w] = c1053obus[data_w*2 +:data_w];
assign c1053ibus[temp_w*3 +:temp_w] = v910obus[temp_w*5 +:temp_w];
assign v910ibus[data_w*5 +:data_w] = c1053obus[data_w*3 +:data_w];
assign c1053ibus[temp_w*4 +:temp_w] = v2205obus[temp_w*1 +:temp_w];
assign v2205ibus[data_w*1 +:data_w] = c1053obus[data_w*4 +:data_w];
assign c1053ibus[temp_w*5 +:temp_w] = v2301obus[temp_w*0 +:temp_w];
assign v2301ibus[data_w*0 +:data_w] = c1053obus[data_w*5 +:data_w];
assign c1054ibus[temp_w*0 +:temp_w] = v197obus[temp_w*5 +:temp_w];
assign v197ibus[data_w*5 +:data_w] = c1054obus[data_w*0 +:data_w];
assign c1054ibus[temp_w*1 +:temp_w] = v351obus[temp_w*2 +:temp_w];
assign v351ibus[data_w*2 +:data_w] = c1054obus[data_w*1 +:data_w];
assign c1054ibus[temp_w*2 +:temp_w] = v805obus[temp_w*2 +:temp_w];
assign v805ibus[data_w*2 +:data_w] = c1054obus[data_w*2 +:data_w];
assign c1054ibus[temp_w*3 +:temp_w] = v911obus[temp_w*5 +:temp_w];
assign v911ibus[data_w*5 +:data_w] = c1054obus[data_w*3 +:data_w];
assign c1054ibus[temp_w*4 +:temp_w] = v2206obus[temp_w*1 +:temp_w];
assign v2206ibus[data_w*1 +:data_w] = c1054obus[data_w*4 +:data_w];
assign c1054ibus[temp_w*5 +:temp_w] = v2302obus[temp_w*0 +:temp_w];
assign v2302ibus[data_w*0 +:data_w] = c1054obus[data_w*5 +:data_w];
assign c1055ibus[temp_w*0 +:temp_w] = v198obus[temp_w*5 +:temp_w];
assign v198ibus[data_w*5 +:data_w] = c1055obus[data_w*0 +:data_w];
assign c1055ibus[temp_w*1 +:temp_w] = v352obus[temp_w*2 +:temp_w];
assign v352ibus[data_w*2 +:data_w] = c1055obus[data_w*1 +:data_w];
assign c1055ibus[temp_w*2 +:temp_w] = v806obus[temp_w*2 +:temp_w];
assign v806ibus[data_w*2 +:data_w] = c1055obus[data_w*2 +:data_w];
assign c1055ibus[temp_w*3 +:temp_w] = v912obus[temp_w*5 +:temp_w];
assign v912ibus[data_w*5 +:data_w] = c1055obus[data_w*3 +:data_w];
assign c1055ibus[temp_w*4 +:temp_w] = v2207obus[temp_w*1 +:temp_w];
assign v2207ibus[data_w*1 +:data_w] = c1055obus[data_w*4 +:data_w];
assign c1055ibus[temp_w*5 +:temp_w] = v2303obus[temp_w*0 +:temp_w];
assign v2303ibus[data_w*0 +:data_w] = c1055obus[data_w*5 +:data_w];
assign c1056ibus[temp_w*0 +:temp_w] = v43obus[temp_w*2 +:temp_w];
assign v43ibus[data_w*2 +:data_w] = c1056obus[data_w*0 +:data_w];
assign c1056ibus[temp_w*1 +:temp_w] = v546obus[temp_w*5 +:temp_w];
assign v546ibus[data_w*5 +:data_w] = c1056obus[data_w*1 +:data_w];
assign c1056ibus[temp_w*2 +:temp_w] = v713obus[temp_w*5 +:temp_w];
assign v713ibus[data_w*5 +:data_w] = c1056obus[data_w*2 +:data_w];
assign c1056ibus[temp_w*3 +:temp_w] = v1082obus[temp_w*5 +:temp_w];
assign v1082ibus[data_w*5 +:data_w] = c1056obus[data_w*3 +:data_w];
assign c1056ibus[temp_w*4 +:temp_w] = v1159obus[temp_w*2 +:temp_w];
assign v1159ibus[data_w*2 +:data_w] = c1056obus[data_w*4 +:data_w];
assign c1056ibus[temp_w*5 +:temp_w] = v2208obus[temp_w*1 +:temp_w];
assign v2208ibus[data_w*1 +:data_w] = c1056obus[data_w*5 +:data_w];
assign c1057ibus[temp_w*0 +:temp_w] = v44obus[temp_w*2 +:temp_w];
assign v44ibus[data_w*2 +:data_w] = c1057obus[data_w*0 +:data_w];
assign c1057ibus[temp_w*1 +:temp_w] = v547obus[temp_w*5 +:temp_w];
assign v547ibus[data_w*5 +:data_w] = c1057obus[data_w*1 +:data_w];
assign c1057ibus[temp_w*2 +:temp_w] = v714obus[temp_w*5 +:temp_w];
assign v714ibus[data_w*5 +:data_w] = c1057obus[data_w*2 +:data_w];
assign c1057ibus[temp_w*3 +:temp_w] = v1083obus[temp_w*5 +:temp_w];
assign v1083ibus[data_w*5 +:data_w] = c1057obus[data_w*3 +:data_w];
assign c1057ibus[temp_w*4 +:temp_w] = v1160obus[temp_w*2 +:temp_w];
assign v1160ibus[data_w*2 +:data_w] = c1057obus[data_w*4 +:data_w];
assign c1057ibus[temp_w*5 +:temp_w] = v2209obus[temp_w*1 +:temp_w];
assign v2209ibus[data_w*1 +:data_w] = c1057obus[data_w*5 +:data_w];
assign c1058ibus[temp_w*0 +:temp_w] = v45obus[temp_w*2 +:temp_w];
assign v45ibus[data_w*2 +:data_w] = c1058obus[data_w*0 +:data_w];
assign c1058ibus[temp_w*1 +:temp_w] = v548obus[temp_w*5 +:temp_w];
assign v548ibus[data_w*5 +:data_w] = c1058obus[data_w*1 +:data_w];
assign c1058ibus[temp_w*2 +:temp_w] = v715obus[temp_w*5 +:temp_w];
assign v715ibus[data_w*5 +:data_w] = c1058obus[data_w*2 +:data_w];
assign c1058ibus[temp_w*3 +:temp_w] = v1084obus[temp_w*5 +:temp_w];
assign v1084ibus[data_w*5 +:data_w] = c1058obus[data_w*3 +:data_w];
assign c1058ibus[temp_w*4 +:temp_w] = v1161obus[temp_w*2 +:temp_w];
assign v1161ibus[data_w*2 +:data_w] = c1058obus[data_w*4 +:data_w];
assign c1058ibus[temp_w*5 +:temp_w] = v2210obus[temp_w*1 +:temp_w];
assign v2210ibus[data_w*1 +:data_w] = c1058obus[data_w*5 +:data_w];
assign c1059ibus[temp_w*0 +:temp_w] = v46obus[temp_w*2 +:temp_w];
assign v46ibus[data_w*2 +:data_w] = c1059obus[data_w*0 +:data_w];
assign c1059ibus[temp_w*1 +:temp_w] = v549obus[temp_w*5 +:temp_w];
assign v549ibus[data_w*5 +:data_w] = c1059obus[data_w*1 +:data_w];
assign c1059ibus[temp_w*2 +:temp_w] = v716obus[temp_w*5 +:temp_w];
assign v716ibus[data_w*5 +:data_w] = c1059obus[data_w*2 +:data_w];
assign c1059ibus[temp_w*3 +:temp_w] = v1085obus[temp_w*5 +:temp_w];
assign v1085ibus[data_w*5 +:data_w] = c1059obus[data_w*3 +:data_w];
assign c1059ibus[temp_w*4 +:temp_w] = v1162obus[temp_w*2 +:temp_w];
assign v1162ibus[data_w*2 +:data_w] = c1059obus[data_w*4 +:data_w];
assign c1059ibus[temp_w*5 +:temp_w] = v2211obus[temp_w*1 +:temp_w];
assign v2211ibus[data_w*1 +:data_w] = c1059obus[data_w*5 +:data_w];
assign c1060ibus[temp_w*0 +:temp_w] = v47obus[temp_w*2 +:temp_w];
assign v47ibus[data_w*2 +:data_w] = c1060obus[data_w*0 +:data_w];
assign c1060ibus[temp_w*1 +:temp_w] = v550obus[temp_w*5 +:temp_w];
assign v550ibus[data_w*5 +:data_w] = c1060obus[data_w*1 +:data_w];
assign c1060ibus[temp_w*2 +:temp_w] = v717obus[temp_w*5 +:temp_w];
assign v717ibus[data_w*5 +:data_w] = c1060obus[data_w*2 +:data_w];
assign c1060ibus[temp_w*3 +:temp_w] = v1086obus[temp_w*5 +:temp_w];
assign v1086ibus[data_w*5 +:data_w] = c1060obus[data_w*3 +:data_w];
assign c1060ibus[temp_w*4 +:temp_w] = v1163obus[temp_w*2 +:temp_w];
assign v1163ibus[data_w*2 +:data_w] = c1060obus[data_w*4 +:data_w];
assign c1060ibus[temp_w*5 +:temp_w] = v2212obus[temp_w*1 +:temp_w];
assign v2212ibus[data_w*1 +:data_w] = c1060obus[data_w*5 +:data_w];
assign c1061ibus[temp_w*0 +:temp_w] = v48obus[temp_w*2 +:temp_w];
assign v48ibus[data_w*2 +:data_w] = c1061obus[data_w*0 +:data_w];
assign c1061ibus[temp_w*1 +:temp_w] = v551obus[temp_w*5 +:temp_w];
assign v551ibus[data_w*5 +:data_w] = c1061obus[data_w*1 +:data_w];
assign c1061ibus[temp_w*2 +:temp_w] = v718obus[temp_w*5 +:temp_w];
assign v718ibus[data_w*5 +:data_w] = c1061obus[data_w*2 +:data_w];
assign c1061ibus[temp_w*3 +:temp_w] = v1087obus[temp_w*5 +:temp_w];
assign v1087ibus[data_w*5 +:data_w] = c1061obus[data_w*3 +:data_w];
assign c1061ibus[temp_w*4 +:temp_w] = v1164obus[temp_w*2 +:temp_w];
assign v1164ibus[data_w*2 +:data_w] = c1061obus[data_w*4 +:data_w];
assign c1061ibus[temp_w*5 +:temp_w] = v2213obus[temp_w*1 +:temp_w];
assign v2213ibus[data_w*1 +:data_w] = c1061obus[data_w*5 +:data_w];
assign c1062ibus[temp_w*0 +:temp_w] = v49obus[temp_w*2 +:temp_w];
assign v49ibus[data_w*2 +:data_w] = c1062obus[data_w*0 +:data_w];
assign c1062ibus[temp_w*1 +:temp_w] = v552obus[temp_w*5 +:temp_w];
assign v552ibus[data_w*5 +:data_w] = c1062obus[data_w*1 +:data_w];
assign c1062ibus[temp_w*2 +:temp_w] = v719obus[temp_w*5 +:temp_w];
assign v719ibus[data_w*5 +:data_w] = c1062obus[data_w*2 +:data_w];
assign c1062ibus[temp_w*3 +:temp_w] = v1088obus[temp_w*5 +:temp_w];
assign v1088ibus[data_w*5 +:data_w] = c1062obus[data_w*3 +:data_w];
assign c1062ibus[temp_w*4 +:temp_w] = v1165obus[temp_w*2 +:temp_w];
assign v1165ibus[data_w*2 +:data_w] = c1062obus[data_w*4 +:data_w];
assign c1062ibus[temp_w*5 +:temp_w] = v2214obus[temp_w*1 +:temp_w];
assign v2214ibus[data_w*1 +:data_w] = c1062obus[data_w*5 +:data_w];
assign c1063ibus[temp_w*0 +:temp_w] = v50obus[temp_w*2 +:temp_w];
assign v50ibus[data_w*2 +:data_w] = c1063obus[data_w*0 +:data_w];
assign c1063ibus[temp_w*1 +:temp_w] = v553obus[temp_w*5 +:temp_w];
assign v553ibus[data_w*5 +:data_w] = c1063obus[data_w*1 +:data_w];
assign c1063ibus[temp_w*2 +:temp_w] = v720obus[temp_w*5 +:temp_w];
assign v720ibus[data_w*5 +:data_w] = c1063obus[data_w*2 +:data_w];
assign c1063ibus[temp_w*3 +:temp_w] = v1089obus[temp_w*5 +:temp_w];
assign v1089ibus[data_w*5 +:data_w] = c1063obus[data_w*3 +:data_w];
assign c1063ibus[temp_w*4 +:temp_w] = v1166obus[temp_w*2 +:temp_w];
assign v1166ibus[data_w*2 +:data_w] = c1063obus[data_w*4 +:data_w];
assign c1063ibus[temp_w*5 +:temp_w] = v2215obus[temp_w*1 +:temp_w];
assign v2215ibus[data_w*1 +:data_w] = c1063obus[data_w*5 +:data_w];
assign c1064ibus[temp_w*0 +:temp_w] = v51obus[temp_w*2 +:temp_w];
assign v51ibus[data_w*2 +:data_w] = c1064obus[data_w*0 +:data_w];
assign c1064ibus[temp_w*1 +:temp_w] = v554obus[temp_w*5 +:temp_w];
assign v554ibus[data_w*5 +:data_w] = c1064obus[data_w*1 +:data_w];
assign c1064ibus[temp_w*2 +:temp_w] = v721obus[temp_w*5 +:temp_w];
assign v721ibus[data_w*5 +:data_w] = c1064obus[data_w*2 +:data_w];
assign c1064ibus[temp_w*3 +:temp_w] = v1090obus[temp_w*5 +:temp_w];
assign v1090ibus[data_w*5 +:data_w] = c1064obus[data_w*3 +:data_w];
assign c1064ibus[temp_w*4 +:temp_w] = v1167obus[temp_w*2 +:temp_w];
assign v1167ibus[data_w*2 +:data_w] = c1064obus[data_w*4 +:data_w];
assign c1064ibus[temp_w*5 +:temp_w] = v2216obus[temp_w*1 +:temp_w];
assign v2216ibus[data_w*1 +:data_w] = c1064obus[data_w*5 +:data_w];
assign c1065ibus[temp_w*0 +:temp_w] = v52obus[temp_w*2 +:temp_w];
assign v52ibus[data_w*2 +:data_w] = c1065obus[data_w*0 +:data_w];
assign c1065ibus[temp_w*1 +:temp_w] = v555obus[temp_w*5 +:temp_w];
assign v555ibus[data_w*5 +:data_w] = c1065obus[data_w*1 +:data_w];
assign c1065ibus[temp_w*2 +:temp_w] = v722obus[temp_w*5 +:temp_w];
assign v722ibus[data_w*5 +:data_w] = c1065obus[data_w*2 +:data_w];
assign c1065ibus[temp_w*3 +:temp_w] = v1091obus[temp_w*5 +:temp_w];
assign v1091ibus[data_w*5 +:data_w] = c1065obus[data_w*3 +:data_w];
assign c1065ibus[temp_w*4 +:temp_w] = v1168obus[temp_w*2 +:temp_w];
assign v1168ibus[data_w*2 +:data_w] = c1065obus[data_w*4 +:data_w];
assign c1065ibus[temp_w*5 +:temp_w] = v2217obus[temp_w*1 +:temp_w];
assign v2217ibus[data_w*1 +:data_w] = c1065obus[data_w*5 +:data_w];
assign c1066ibus[temp_w*0 +:temp_w] = v53obus[temp_w*2 +:temp_w];
assign v53ibus[data_w*2 +:data_w] = c1066obus[data_w*0 +:data_w];
assign c1066ibus[temp_w*1 +:temp_w] = v556obus[temp_w*5 +:temp_w];
assign v556ibus[data_w*5 +:data_w] = c1066obus[data_w*1 +:data_w];
assign c1066ibus[temp_w*2 +:temp_w] = v723obus[temp_w*5 +:temp_w];
assign v723ibus[data_w*5 +:data_w] = c1066obus[data_w*2 +:data_w];
assign c1066ibus[temp_w*3 +:temp_w] = v1092obus[temp_w*5 +:temp_w];
assign v1092ibus[data_w*5 +:data_w] = c1066obus[data_w*3 +:data_w];
assign c1066ibus[temp_w*4 +:temp_w] = v1169obus[temp_w*2 +:temp_w];
assign v1169ibus[data_w*2 +:data_w] = c1066obus[data_w*4 +:data_w];
assign c1066ibus[temp_w*5 +:temp_w] = v2218obus[temp_w*1 +:temp_w];
assign v2218ibus[data_w*1 +:data_w] = c1066obus[data_w*5 +:data_w];
assign c1067ibus[temp_w*0 +:temp_w] = v54obus[temp_w*2 +:temp_w];
assign v54ibus[data_w*2 +:data_w] = c1067obus[data_w*0 +:data_w];
assign c1067ibus[temp_w*1 +:temp_w] = v557obus[temp_w*5 +:temp_w];
assign v557ibus[data_w*5 +:data_w] = c1067obus[data_w*1 +:data_w];
assign c1067ibus[temp_w*2 +:temp_w] = v724obus[temp_w*5 +:temp_w];
assign v724ibus[data_w*5 +:data_w] = c1067obus[data_w*2 +:data_w];
assign c1067ibus[temp_w*3 +:temp_w] = v1093obus[temp_w*5 +:temp_w];
assign v1093ibus[data_w*5 +:data_w] = c1067obus[data_w*3 +:data_w];
assign c1067ibus[temp_w*4 +:temp_w] = v1170obus[temp_w*2 +:temp_w];
assign v1170ibus[data_w*2 +:data_w] = c1067obus[data_w*4 +:data_w];
assign c1067ibus[temp_w*5 +:temp_w] = v2219obus[temp_w*1 +:temp_w];
assign v2219ibus[data_w*1 +:data_w] = c1067obus[data_w*5 +:data_w];
assign c1068ibus[temp_w*0 +:temp_w] = v55obus[temp_w*2 +:temp_w];
assign v55ibus[data_w*2 +:data_w] = c1068obus[data_w*0 +:data_w];
assign c1068ibus[temp_w*1 +:temp_w] = v558obus[temp_w*5 +:temp_w];
assign v558ibus[data_w*5 +:data_w] = c1068obus[data_w*1 +:data_w];
assign c1068ibus[temp_w*2 +:temp_w] = v725obus[temp_w*5 +:temp_w];
assign v725ibus[data_w*5 +:data_w] = c1068obus[data_w*2 +:data_w];
assign c1068ibus[temp_w*3 +:temp_w] = v1094obus[temp_w*5 +:temp_w];
assign v1094ibus[data_w*5 +:data_w] = c1068obus[data_w*3 +:data_w];
assign c1068ibus[temp_w*4 +:temp_w] = v1171obus[temp_w*2 +:temp_w];
assign v1171ibus[data_w*2 +:data_w] = c1068obus[data_w*4 +:data_w];
assign c1068ibus[temp_w*5 +:temp_w] = v2220obus[temp_w*1 +:temp_w];
assign v2220ibus[data_w*1 +:data_w] = c1068obus[data_w*5 +:data_w];
assign c1069ibus[temp_w*0 +:temp_w] = v56obus[temp_w*2 +:temp_w];
assign v56ibus[data_w*2 +:data_w] = c1069obus[data_w*0 +:data_w];
assign c1069ibus[temp_w*1 +:temp_w] = v559obus[temp_w*5 +:temp_w];
assign v559ibus[data_w*5 +:data_w] = c1069obus[data_w*1 +:data_w];
assign c1069ibus[temp_w*2 +:temp_w] = v726obus[temp_w*5 +:temp_w];
assign v726ibus[data_w*5 +:data_w] = c1069obus[data_w*2 +:data_w];
assign c1069ibus[temp_w*3 +:temp_w] = v1095obus[temp_w*5 +:temp_w];
assign v1095ibus[data_w*5 +:data_w] = c1069obus[data_w*3 +:data_w];
assign c1069ibus[temp_w*4 +:temp_w] = v1172obus[temp_w*2 +:temp_w];
assign v1172ibus[data_w*2 +:data_w] = c1069obus[data_w*4 +:data_w];
assign c1069ibus[temp_w*5 +:temp_w] = v2221obus[temp_w*1 +:temp_w];
assign v2221ibus[data_w*1 +:data_w] = c1069obus[data_w*5 +:data_w];
assign c1070ibus[temp_w*0 +:temp_w] = v57obus[temp_w*2 +:temp_w];
assign v57ibus[data_w*2 +:data_w] = c1070obus[data_w*0 +:data_w];
assign c1070ibus[temp_w*1 +:temp_w] = v560obus[temp_w*5 +:temp_w];
assign v560ibus[data_w*5 +:data_w] = c1070obus[data_w*1 +:data_w];
assign c1070ibus[temp_w*2 +:temp_w] = v727obus[temp_w*5 +:temp_w];
assign v727ibus[data_w*5 +:data_w] = c1070obus[data_w*2 +:data_w];
assign c1070ibus[temp_w*3 +:temp_w] = v1096obus[temp_w*5 +:temp_w];
assign v1096ibus[data_w*5 +:data_w] = c1070obus[data_w*3 +:data_w];
assign c1070ibus[temp_w*4 +:temp_w] = v1173obus[temp_w*2 +:temp_w];
assign v1173ibus[data_w*2 +:data_w] = c1070obus[data_w*4 +:data_w];
assign c1070ibus[temp_w*5 +:temp_w] = v2222obus[temp_w*1 +:temp_w];
assign v2222ibus[data_w*1 +:data_w] = c1070obus[data_w*5 +:data_w];
assign c1071ibus[temp_w*0 +:temp_w] = v58obus[temp_w*2 +:temp_w];
assign v58ibus[data_w*2 +:data_w] = c1071obus[data_w*0 +:data_w];
assign c1071ibus[temp_w*1 +:temp_w] = v561obus[temp_w*5 +:temp_w];
assign v561ibus[data_w*5 +:data_w] = c1071obus[data_w*1 +:data_w];
assign c1071ibus[temp_w*2 +:temp_w] = v728obus[temp_w*5 +:temp_w];
assign v728ibus[data_w*5 +:data_w] = c1071obus[data_w*2 +:data_w];
assign c1071ibus[temp_w*3 +:temp_w] = v1097obus[temp_w*5 +:temp_w];
assign v1097ibus[data_w*5 +:data_w] = c1071obus[data_w*3 +:data_w];
assign c1071ibus[temp_w*4 +:temp_w] = v1174obus[temp_w*2 +:temp_w];
assign v1174ibus[data_w*2 +:data_w] = c1071obus[data_w*4 +:data_w];
assign c1071ibus[temp_w*5 +:temp_w] = v2223obus[temp_w*1 +:temp_w];
assign v2223ibus[data_w*1 +:data_w] = c1071obus[data_w*5 +:data_w];
assign c1072ibus[temp_w*0 +:temp_w] = v59obus[temp_w*2 +:temp_w];
assign v59ibus[data_w*2 +:data_w] = c1072obus[data_w*0 +:data_w];
assign c1072ibus[temp_w*1 +:temp_w] = v562obus[temp_w*5 +:temp_w];
assign v562ibus[data_w*5 +:data_w] = c1072obus[data_w*1 +:data_w];
assign c1072ibus[temp_w*2 +:temp_w] = v729obus[temp_w*5 +:temp_w];
assign v729ibus[data_w*5 +:data_w] = c1072obus[data_w*2 +:data_w];
assign c1072ibus[temp_w*3 +:temp_w] = v1098obus[temp_w*5 +:temp_w];
assign v1098ibus[data_w*5 +:data_w] = c1072obus[data_w*3 +:data_w];
assign c1072ibus[temp_w*4 +:temp_w] = v1175obus[temp_w*2 +:temp_w];
assign v1175ibus[data_w*2 +:data_w] = c1072obus[data_w*4 +:data_w];
assign c1072ibus[temp_w*5 +:temp_w] = v2224obus[temp_w*1 +:temp_w];
assign v2224ibus[data_w*1 +:data_w] = c1072obus[data_w*5 +:data_w];
assign c1073ibus[temp_w*0 +:temp_w] = v60obus[temp_w*2 +:temp_w];
assign v60ibus[data_w*2 +:data_w] = c1073obus[data_w*0 +:data_w];
assign c1073ibus[temp_w*1 +:temp_w] = v563obus[temp_w*5 +:temp_w];
assign v563ibus[data_w*5 +:data_w] = c1073obus[data_w*1 +:data_w];
assign c1073ibus[temp_w*2 +:temp_w] = v730obus[temp_w*5 +:temp_w];
assign v730ibus[data_w*5 +:data_w] = c1073obus[data_w*2 +:data_w];
assign c1073ibus[temp_w*3 +:temp_w] = v1099obus[temp_w*5 +:temp_w];
assign v1099ibus[data_w*5 +:data_w] = c1073obus[data_w*3 +:data_w];
assign c1073ibus[temp_w*4 +:temp_w] = v1176obus[temp_w*2 +:temp_w];
assign v1176ibus[data_w*2 +:data_w] = c1073obus[data_w*4 +:data_w];
assign c1073ibus[temp_w*5 +:temp_w] = v2225obus[temp_w*1 +:temp_w];
assign v2225ibus[data_w*1 +:data_w] = c1073obus[data_w*5 +:data_w];
assign c1074ibus[temp_w*0 +:temp_w] = v61obus[temp_w*2 +:temp_w];
assign v61ibus[data_w*2 +:data_w] = c1074obus[data_w*0 +:data_w];
assign c1074ibus[temp_w*1 +:temp_w] = v564obus[temp_w*5 +:temp_w];
assign v564ibus[data_w*5 +:data_w] = c1074obus[data_w*1 +:data_w];
assign c1074ibus[temp_w*2 +:temp_w] = v731obus[temp_w*5 +:temp_w];
assign v731ibus[data_w*5 +:data_w] = c1074obus[data_w*2 +:data_w];
assign c1074ibus[temp_w*3 +:temp_w] = v1100obus[temp_w*5 +:temp_w];
assign v1100ibus[data_w*5 +:data_w] = c1074obus[data_w*3 +:data_w];
assign c1074ibus[temp_w*4 +:temp_w] = v1177obus[temp_w*2 +:temp_w];
assign v1177ibus[data_w*2 +:data_w] = c1074obus[data_w*4 +:data_w];
assign c1074ibus[temp_w*5 +:temp_w] = v2226obus[temp_w*1 +:temp_w];
assign v2226ibus[data_w*1 +:data_w] = c1074obus[data_w*5 +:data_w];
assign c1075ibus[temp_w*0 +:temp_w] = v62obus[temp_w*2 +:temp_w];
assign v62ibus[data_w*2 +:data_w] = c1075obus[data_w*0 +:data_w];
assign c1075ibus[temp_w*1 +:temp_w] = v565obus[temp_w*5 +:temp_w];
assign v565ibus[data_w*5 +:data_w] = c1075obus[data_w*1 +:data_w];
assign c1075ibus[temp_w*2 +:temp_w] = v732obus[temp_w*5 +:temp_w];
assign v732ibus[data_w*5 +:data_w] = c1075obus[data_w*2 +:data_w];
assign c1075ibus[temp_w*3 +:temp_w] = v1101obus[temp_w*5 +:temp_w];
assign v1101ibus[data_w*5 +:data_w] = c1075obus[data_w*3 +:data_w];
assign c1075ibus[temp_w*4 +:temp_w] = v1178obus[temp_w*2 +:temp_w];
assign v1178ibus[data_w*2 +:data_w] = c1075obus[data_w*4 +:data_w];
assign c1075ibus[temp_w*5 +:temp_w] = v2227obus[temp_w*1 +:temp_w];
assign v2227ibus[data_w*1 +:data_w] = c1075obus[data_w*5 +:data_w];
assign c1076ibus[temp_w*0 +:temp_w] = v63obus[temp_w*2 +:temp_w];
assign v63ibus[data_w*2 +:data_w] = c1076obus[data_w*0 +:data_w];
assign c1076ibus[temp_w*1 +:temp_w] = v566obus[temp_w*5 +:temp_w];
assign v566ibus[data_w*5 +:data_w] = c1076obus[data_w*1 +:data_w];
assign c1076ibus[temp_w*2 +:temp_w] = v733obus[temp_w*5 +:temp_w];
assign v733ibus[data_w*5 +:data_w] = c1076obus[data_w*2 +:data_w];
assign c1076ibus[temp_w*3 +:temp_w] = v1102obus[temp_w*5 +:temp_w];
assign v1102ibus[data_w*5 +:data_w] = c1076obus[data_w*3 +:data_w];
assign c1076ibus[temp_w*4 +:temp_w] = v1179obus[temp_w*2 +:temp_w];
assign v1179ibus[data_w*2 +:data_w] = c1076obus[data_w*4 +:data_w];
assign c1076ibus[temp_w*5 +:temp_w] = v2228obus[temp_w*1 +:temp_w];
assign v2228ibus[data_w*1 +:data_w] = c1076obus[data_w*5 +:data_w];
assign c1077ibus[temp_w*0 +:temp_w] = v64obus[temp_w*2 +:temp_w];
assign v64ibus[data_w*2 +:data_w] = c1077obus[data_w*0 +:data_w];
assign c1077ibus[temp_w*1 +:temp_w] = v567obus[temp_w*5 +:temp_w];
assign v567ibus[data_w*5 +:data_w] = c1077obus[data_w*1 +:data_w];
assign c1077ibus[temp_w*2 +:temp_w] = v734obus[temp_w*5 +:temp_w];
assign v734ibus[data_w*5 +:data_w] = c1077obus[data_w*2 +:data_w];
assign c1077ibus[temp_w*3 +:temp_w] = v1103obus[temp_w*5 +:temp_w];
assign v1103ibus[data_w*5 +:data_w] = c1077obus[data_w*3 +:data_w];
assign c1077ibus[temp_w*4 +:temp_w] = v1180obus[temp_w*2 +:temp_w];
assign v1180ibus[data_w*2 +:data_w] = c1077obus[data_w*4 +:data_w];
assign c1077ibus[temp_w*5 +:temp_w] = v2229obus[temp_w*1 +:temp_w];
assign v2229ibus[data_w*1 +:data_w] = c1077obus[data_w*5 +:data_w];
assign c1078ibus[temp_w*0 +:temp_w] = v65obus[temp_w*2 +:temp_w];
assign v65ibus[data_w*2 +:data_w] = c1078obus[data_w*0 +:data_w];
assign c1078ibus[temp_w*1 +:temp_w] = v568obus[temp_w*5 +:temp_w];
assign v568ibus[data_w*5 +:data_w] = c1078obus[data_w*1 +:data_w];
assign c1078ibus[temp_w*2 +:temp_w] = v735obus[temp_w*5 +:temp_w];
assign v735ibus[data_w*5 +:data_w] = c1078obus[data_w*2 +:data_w];
assign c1078ibus[temp_w*3 +:temp_w] = v1104obus[temp_w*5 +:temp_w];
assign v1104ibus[data_w*5 +:data_w] = c1078obus[data_w*3 +:data_w];
assign c1078ibus[temp_w*4 +:temp_w] = v1181obus[temp_w*2 +:temp_w];
assign v1181ibus[data_w*2 +:data_w] = c1078obus[data_w*4 +:data_w];
assign c1078ibus[temp_w*5 +:temp_w] = v2230obus[temp_w*1 +:temp_w];
assign v2230ibus[data_w*1 +:data_w] = c1078obus[data_w*5 +:data_w];
assign c1079ibus[temp_w*0 +:temp_w] = v66obus[temp_w*2 +:temp_w];
assign v66ibus[data_w*2 +:data_w] = c1079obus[data_w*0 +:data_w];
assign c1079ibus[temp_w*1 +:temp_w] = v569obus[temp_w*5 +:temp_w];
assign v569ibus[data_w*5 +:data_w] = c1079obus[data_w*1 +:data_w];
assign c1079ibus[temp_w*2 +:temp_w] = v736obus[temp_w*5 +:temp_w];
assign v736ibus[data_w*5 +:data_w] = c1079obus[data_w*2 +:data_w];
assign c1079ibus[temp_w*3 +:temp_w] = v1105obus[temp_w*5 +:temp_w];
assign v1105ibus[data_w*5 +:data_w] = c1079obus[data_w*3 +:data_w];
assign c1079ibus[temp_w*4 +:temp_w] = v1182obus[temp_w*2 +:temp_w];
assign v1182ibus[data_w*2 +:data_w] = c1079obus[data_w*4 +:data_w];
assign c1079ibus[temp_w*5 +:temp_w] = v2231obus[temp_w*1 +:temp_w];
assign v2231ibus[data_w*1 +:data_w] = c1079obus[data_w*5 +:data_w];
assign c1080ibus[temp_w*0 +:temp_w] = v67obus[temp_w*2 +:temp_w];
assign v67ibus[data_w*2 +:data_w] = c1080obus[data_w*0 +:data_w];
assign c1080ibus[temp_w*1 +:temp_w] = v570obus[temp_w*5 +:temp_w];
assign v570ibus[data_w*5 +:data_w] = c1080obus[data_w*1 +:data_w];
assign c1080ibus[temp_w*2 +:temp_w] = v737obus[temp_w*5 +:temp_w];
assign v737ibus[data_w*5 +:data_w] = c1080obus[data_w*2 +:data_w];
assign c1080ibus[temp_w*3 +:temp_w] = v1106obus[temp_w*5 +:temp_w];
assign v1106ibus[data_w*5 +:data_w] = c1080obus[data_w*3 +:data_w];
assign c1080ibus[temp_w*4 +:temp_w] = v1183obus[temp_w*2 +:temp_w];
assign v1183ibus[data_w*2 +:data_w] = c1080obus[data_w*4 +:data_w];
assign c1080ibus[temp_w*5 +:temp_w] = v2232obus[temp_w*1 +:temp_w];
assign v2232ibus[data_w*1 +:data_w] = c1080obus[data_w*5 +:data_w];
assign c1081ibus[temp_w*0 +:temp_w] = v68obus[temp_w*2 +:temp_w];
assign v68ibus[data_w*2 +:data_w] = c1081obus[data_w*0 +:data_w];
assign c1081ibus[temp_w*1 +:temp_w] = v571obus[temp_w*5 +:temp_w];
assign v571ibus[data_w*5 +:data_w] = c1081obus[data_w*1 +:data_w];
assign c1081ibus[temp_w*2 +:temp_w] = v738obus[temp_w*5 +:temp_w];
assign v738ibus[data_w*5 +:data_w] = c1081obus[data_w*2 +:data_w];
assign c1081ibus[temp_w*3 +:temp_w] = v1107obus[temp_w*5 +:temp_w];
assign v1107ibus[data_w*5 +:data_w] = c1081obus[data_w*3 +:data_w];
assign c1081ibus[temp_w*4 +:temp_w] = v1184obus[temp_w*2 +:temp_w];
assign v1184ibus[data_w*2 +:data_w] = c1081obus[data_w*4 +:data_w];
assign c1081ibus[temp_w*5 +:temp_w] = v2233obus[temp_w*1 +:temp_w];
assign v2233ibus[data_w*1 +:data_w] = c1081obus[data_w*5 +:data_w];
assign c1082ibus[temp_w*0 +:temp_w] = v69obus[temp_w*2 +:temp_w];
assign v69ibus[data_w*2 +:data_w] = c1082obus[data_w*0 +:data_w];
assign c1082ibus[temp_w*1 +:temp_w] = v572obus[temp_w*5 +:temp_w];
assign v572ibus[data_w*5 +:data_w] = c1082obus[data_w*1 +:data_w];
assign c1082ibus[temp_w*2 +:temp_w] = v739obus[temp_w*5 +:temp_w];
assign v739ibus[data_w*5 +:data_w] = c1082obus[data_w*2 +:data_w];
assign c1082ibus[temp_w*3 +:temp_w] = v1108obus[temp_w*5 +:temp_w];
assign v1108ibus[data_w*5 +:data_w] = c1082obus[data_w*3 +:data_w];
assign c1082ibus[temp_w*4 +:temp_w] = v1185obus[temp_w*2 +:temp_w];
assign v1185ibus[data_w*2 +:data_w] = c1082obus[data_w*4 +:data_w];
assign c1082ibus[temp_w*5 +:temp_w] = v2234obus[temp_w*1 +:temp_w];
assign v2234ibus[data_w*1 +:data_w] = c1082obus[data_w*5 +:data_w];
assign c1083ibus[temp_w*0 +:temp_w] = v70obus[temp_w*2 +:temp_w];
assign v70ibus[data_w*2 +:data_w] = c1083obus[data_w*0 +:data_w];
assign c1083ibus[temp_w*1 +:temp_w] = v573obus[temp_w*5 +:temp_w];
assign v573ibus[data_w*5 +:data_w] = c1083obus[data_w*1 +:data_w];
assign c1083ibus[temp_w*2 +:temp_w] = v740obus[temp_w*5 +:temp_w];
assign v740ibus[data_w*5 +:data_w] = c1083obus[data_w*2 +:data_w];
assign c1083ibus[temp_w*3 +:temp_w] = v1109obus[temp_w*5 +:temp_w];
assign v1109ibus[data_w*5 +:data_w] = c1083obus[data_w*3 +:data_w];
assign c1083ibus[temp_w*4 +:temp_w] = v1186obus[temp_w*2 +:temp_w];
assign v1186ibus[data_w*2 +:data_w] = c1083obus[data_w*4 +:data_w];
assign c1083ibus[temp_w*5 +:temp_w] = v2235obus[temp_w*1 +:temp_w];
assign v2235ibus[data_w*1 +:data_w] = c1083obus[data_w*5 +:data_w];
assign c1084ibus[temp_w*0 +:temp_w] = v71obus[temp_w*2 +:temp_w];
assign v71ibus[data_w*2 +:data_w] = c1084obus[data_w*0 +:data_w];
assign c1084ibus[temp_w*1 +:temp_w] = v574obus[temp_w*5 +:temp_w];
assign v574ibus[data_w*5 +:data_w] = c1084obus[data_w*1 +:data_w];
assign c1084ibus[temp_w*2 +:temp_w] = v741obus[temp_w*5 +:temp_w];
assign v741ibus[data_w*5 +:data_w] = c1084obus[data_w*2 +:data_w];
assign c1084ibus[temp_w*3 +:temp_w] = v1110obus[temp_w*5 +:temp_w];
assign v1110ibus[data_w*5 +:data_w] = c1084obus[data_w*3 +:data_w];
assign c1084ibus[temp_w*4 +:temp_w] = v1187obus[temp_w*2 +:temp_w];
assign v1187ibus[data_w*2 +:data_w] = c1084obus[data_w*4 +:data_w];
assign c1084ibus[temp_w*5 +:temp_w] = v2236obus[temp_w*1 +:temp_w];
assign v2236ibus[data_w*1 +:data_w] = c1084obus[data_w*5 +:data_w];
assign c1085ibus[temp_w*0 +:temp_w] = v72obus[temp_w*2 +:temp_w];
assign v72ibus[data_w*2 +:data_w] = c1085obus[data_w*0 +:data_w];
assign c1085ibus[temp_w*1 +:temp_w] = v575obus[temp_w*5 +:temp_w];
assign v575ibus[data_w*5 +:data_w] = c1085obus[data_w*1 +:data_w];
assign c1085ibus[temp_w*2 +:temp_w] = v742obus[temp_w*5 +:temp_w];
assign v742ibus[data_w*5 +:data_w] = c1085obus[data_w*2 +:data_w];
assign c1085ibus[temp_w*3 +:temp_w] = v1111obus[temp_w*5 +:temp_w];
assign v1111ibus[data_w*5 +:data_w] = c1085obus[data_w*3 +:data_w];
assign c1085ibus[temp_w*4 +:temp_w] = v1188obus[temp_w*2 +:temp_w];
assign v1188ibus[data_w*2 +:data_w] = c1085obus[data_w*4 +:data_w];
assign c1085ibus[temp_w*5 +:temp_w] = v2237obus[temp_w*1 +:temp_w];
assign v2237ibus[data_w*1 +:data_w] = c1085obus[data_w*5 +:data_w];
assign c1086ibus[temp_w*0 +:temp_w] = v73obus[temp_w*2 +:temp_w];
assign v73ibus[data_w*2 +:data_w] = c1086obus[data_w*0 +:data_w];
assign c1086ibus[temp_w*1 +:temp_w] = v480obus[temp_w*5 +:temp_w];
assign v480ibus[data_w*5 +:data_w] = c1086obus[data_w*1 +:data_w];
assign c1086ibus[temp_w*2 +:temp_w] = v743obus[temp_w*5 +:temp_w];
assign v743ibus[data_w*5 +:data_w] = c1086obus[data_w*2 +:data_w];
assign c1086ibus[temp_w*3 +:temp_w] = v1112obus[temp_w*5 +:temp_w];
assign v1112ibus[data_w*5 +:data_w] = c1086obus[data_w*3 +:data_w];
assign c1086ibus[temp_w*4 +:temp_w] = v1189obus[temp_w*2 +:temp_w];
assign v1189ibus[data_w*2 +:data_w] = c1086obus[data_w*4 +:data_w];
assign c1086ibus[temp_w*5 +:temp_w] = v2238obus[temp_w*1 +:temp_w];
assign v2238ibus[data_w*1 +:data_w] = c1086obus[data_w*5 +:data_w];
assign c1087ibus[temp_w*0 +:temp_w] = v74obus[temp_w*2 +:temp_w];
assign v74ibus[data_w*2 +:data_w] = c1087obus[data_w*0 +:data_w];
assign c1087ibus[temp_w*1 +:temp_w] = v481obus[temp_w*5 +:temp_w];
assign v481ibus[data_w*5 +:data_w] = c1087obus[data_w*1 +:data_w];
assign c1087ibus[temp_w*2 +:temp_w] = v744obus[temp_w*5 +:temp_w];
assign v744ibus[data_w*5 +:data_w] = c1087obus[data_w*2 +:data_w];
assign c1087ibus[temp_w*3 +:temp_w] = v1113obus[temp_w*5 +:temp_w];
assign v1113ibus[data_w*5 +:data_w] = c1087obus[data_w*3 +:data_w];
assign c1087ibus[temp_w*4 +:temp_w] = v1190obus[temp_w*2 +:temp_w];
assign v1190ibus[data_w*2 +:data_w] = c1087obus[data_w*4 +:data_w];
assign c1087ibus[temp_w*5 +:temp_w] = v2239obus[temp_w*1 +:temp_w];
assign v2239ibus[data_w*1 +:data_w] = c1087obus[data_w*5 +:data_w];
assign c1088ibus[temp_w*0 +:temp_w] = v75obus[temp_w*2 +:temp_w];
assign v75ibus[data_w*2 +:data_w] = c1088obus[data_w*0 +:data_w];
assign c1088ibus[temp_w*1 +:temp_w] = v482obus[temp_w*5 +:temp_w];
assign v482ibus[data_w*5 +:data_w] = c1088obus[data_w*1 +:data_w];
assign c1088ibus[temp_w*2 +:temp_w] = v745obus[temp_w*5 +:temp_w];
assign v745ibus[data_w*5 +:data_w] = c1088obus[data_w*2 +:data_w];
assign c1088ibus[temp_w*3 +:temp_w] = v1114obus[temp_w*5 +:temp_w];
assign v1114ibus[data_w*5 +:data_w] = c1088obus[data_w*3 +:data_w];
assign c1088ibus[temp_w*4 +:temp_w] = v1191obus[temp_w*2 +:temp_w];
assign v1191ibus[data_w*2 +:data_w] = c1088obus[data_w*4 +:data_w];
assign c1088ibus[temp_w*5 +:temp_w] = v2240obus[temp_w*1 +:temp_w];
assign v2240ibus[data_w*1 +:data_w] = c1088obus[data_w*5 +:data_w];
assign c1089ibus[temp_w*0 +:temp_w] = v76obus[temp_w*2 +:temp_w];
assign v76ibus[data_w*2 +:data_w] = c1089obus[data_w*0 +:data_w];
assign c1089ibus[temp_w*1 +:temp_w] = v483obus[temp_w*5 +:temp_w];
assign v483ibus[data_w*5 +:data_w] = c1089obus[data_w*1 +:data_w];
assign c1089ibus[temp_w*2 +:temp_w] = v746obus[temp_w*5 +:temp_w];
assign v746ibus[data_w*5 +:data_w] = c1089obus[data_w*2 +:data_w];
assign c1089ibus[temp_w*3 +:temp_w] = v1115obus[temp_w*5 +:temp_w];
assign v1115ibus[data_w*5 +:data_w] = c1089obus[data_w*3 +:data_w];
assign c1089ibus[temp_w*4 +:temp_w] = v1192obus[temp_w*2 +:temp_w];
assign v1192ibus[data_w*2 +:data_w] = c1089obus[data_w*4 +:data_w];
assign c1089ibus[temp_w*5 +:temp_w] = v2241obus[temp_w*1 +:temp_w];
assign v2241ibus[data_w*1 +:data_w] = c1089obus[data_w*5 +:data_w];
assign c1090ibus[temp_w*0 +:temp_w] = v77obus[temp_w*2 +:temp_w];
assign v77ibus[data_w*2 +:data_w] = c1090obus[data_w*0 +:data_w];
assign c1090ibus[temp_w*1 +:temp_w] = v484obus[temp_w*5 +:temp_w];
assign v484ibus[data_w*5 +:data_w] = c1090obus[data_w*1 +:data_w];
assign c1090ibus[temp_w*2 +:temp_w] = v747obus[temp_w*5 +:temp_w];
assign v747ibus[data_w*5 +:data_w] = c1090obus[data_w*2 +:data_w];
assign c1090ibus[temp_w*3 +:temp_w] = v1116obus[temp_w*5 +:temp_w];
assign v1116ibus[data_w*5 +:data_w] = c1090obus[data_w*3 +:data_w];
assign c1090ibus[temp_w*4 +:temp_w] = v1193obus[temp_w*2 +:temp_w];
assign v1193ibus[data_w*2 +:data_w] = c1090obus[data_w*4 +:data_w];
assign c1090ibus[temp_w*5 +:temp_w] = v2242obus[temp_w*1 +:temp_w];
assign v2242ibus[data_w*1 +:data_w] = c1090obus[data_w*5 +:data_w];
assign c1091ibus[temp_w*0 +:temp_w] = v78obus[temp_w*2 +:temp_w];
assign v78ibus[data_w*2 +:data_w] = c1091obus[data_w*0 +:data_w];
assign c1091ibus[temp_w*1 +:temp_w] = v485obus[temp_w*5 +:temp_w];
assign v485ibus[data_w*5 +:data_w] = c1091obus[data_w*1 +:data_w];
assign c1091ibus[temp_w*2 +:temp_w] = v748obus[temp_w*5 +:temp_w];
assign v748ibus[data_w*5 +:data_w] = c1091obus[data_w*2 +:data_w];
assign c1091ibus[temp_w*3 +:temp_w] = v1117obus[temp_w*5 +:temp_w];
assign v1117ibus[data_w*5 +:data_w] = c1091obus[data_w*3 +:data_w];
assign c1091ibus[temp_w*4 +:temp_w] = v1194obus[temp_w*2 +:temp_w];
assign v1194ibus[data_w*2 +:data_w] = c1091obus[data_w*4 +:data_w];
assign c1091ibus[temp_w*5 +:temp_w] = v2243obus[temp_w*1 +:temp_w];
assign v2243ibus[data_w*1 +:data_w] = c1091obus[data_w*5 +:data_w];
assign c1092ibus[temp_w*0 +:temp_w] = v79obus[temp_w*2 +:temp_w];
assign v79ibus[data_w*2 +:data_w] = c1092obus[data_w*0 +:data_w];
assign c1092ibus[temp_w*1 +:temp_w] = v486obus[temp_w*5 +:temp_w];
assign v486ibus[data_w*5 +:data_w] = c1092obus[data_w*1 +:data_w];
assign c1092ibus[temp_w*2 +:temp_w] = v749obus[temp_w*5 +:temp_w];
assign v749ibus[data_w*5 +:data_w] = c1092obus[data_w*2 +:data_w];
assign c1092ibus[temp_w*3 +:temp_w] = v1118obus[temp_w*5 +:temp_w];
assign v1118ibus[data_w*5 +:data_w] = c1092obus[data_w*3 +:data_w];
assign c1092ibus[temp_w*4 +:temp_w] = v1195obus[temp_w*2 +:temp_w];
assign v1195ibus[data_w*2 +:data_w] = c1092obus[data_w*4 +:data_w];
assign c1092ibus[temp_w*5 +:temp_w] = v2244obus[temp_w*1 +:temp_w];
assign v2244ibus[data_w*1 +:data_w] = c1092obus[data_w*5 +:data_w];
assign c1093ibus[temp_w*0 +:temp_w] = v80obus[temp_w*2 +:temp_w];
assign v80ibus[data_w*2 +:data_w] = c1093obus[data_w*0 +:data_w];
assign c1093ibus[temp_w*1 +:temp_w] = v487obus[temp_w*5 +:temp_w];
assign v487ibus[data_w*5 +:data_w] = c1093obus[data_w*1 +:data_w];
assign c1093ibus[temp_w*2 +:temp_w] = v750obus[temp_w*5 +:temp_w];
assign v750ibus[data_w*5 +:data_w] = c1093obus[data_w*2 +:data_w];
assign c1093ibus[temp_w*3 +:temp_w] = v1119obus[temp_w*5 +:temp_w];
assign v1119ibus[data_w*5 +:data_w] = c1093obus[data_w*3 +:data_w];
assign c1093ibus[temp_w*4 +:temp_w] = v1196obus[temp_w*2 +:temp_w];
assign v1196ibus[data_w*2 +:data_w] = c1093obus[data_w*4 +:data_w];
assign c1093ibus[temp_w*5 +:temp_w] = v2245obus[temp_w*1 +:temp_w];
assign v2245ibus[data_w*1 +:data_w] = c1093obus[data_w*5 +:data_w];
assign c1094ibus[temp_w*0 +:temp_w] = v81obus[temp_w*2 +:temp_w];
assign v81ibus[data_w*2 +:data_w] = c1094obus[data_w*0 +:data_w];
assign c1094ibus[temp_w*1 +:temp_w] = v488obus[temp_w*5 +:temp_w];
assign v488ibus[data_w*5 +:data_w] = c1094obus[data_w*1 +:data_w];
assign c1094ibus[temp_w*2 +:temp_w] = v751obus[temp_w*5 +:temp_w];
assign v751ibus[data_w*5 +:data_w] = c1094obus[data_w*2 +:data_w];
assign c1094ibus[temp_w*3 +:temp_w] = v1120obus[temp_w*5 +:temp_w];
assign v1120ibus[data_w*5 +:data_w] = c1094obus[data_w*3 +:data_w];
assign c1094ibus[temp_w*4 +:temp_w] = v1197obus[temp_w*2 +:temp_w];
assign v1197ibus[data_w*2 +:data_w] = c1094obus[data_w*4 +:data_w];
assign c1094ibus[temp_w*5 +:temp_w] = v2246obus[temp_w*1 +:temp_w];
assign v2246ibus[data_w*1 +:data_w] = c1094obus[data_w*5 +:data_w];
assign c1095ibus[temp_w*0 +:temp_w] = v82obus[temp_w*2 +:temp_w];
assign v82ibus[data_w*2 +:data_w] = c1095obus[data_w*0 +:data_w];
assign c1095ibus[temp_w*1 +:temp_w] = v489obus[temp_w*5 +:temp_w];
assign v489ibus[data_w*5 +:data_w] = c1095obus[data_w*1 +:data_w];
assign c1095ibus[temp_w*2 +:temp_w] = v752obus[temp_w*5 +:temp_w];
assign v752ibus[data_w*5 +:data_w] = c1095obus[data_w*2 +:data_w];
assign c1095ibus[temp_w*3 +:temp_w] = v1121obus[temp_w*5 +:temp_w];
assign v1121ibus[data_w*5 +:data_w] = c1095obus[data_w*3 +:data_w];
assign c1095ibus[temp_w*4 +:temp_w] = v1198obus[temp_w*2 +:temp_w];
assign v1198ibus[data_w*2 +:data_w] = c1095obus[data_w*4 +:data_w];
assign c1095ibus[temp_w*5 +:temp_w] = v2247obus[temp_w*1 +:temp_w];
assign v2247ibus[data_w*1 +:data_w] = c1095obus[data_w*5 +:data_w];
assign c1096ibus[temp_w*0 +:temp_w] = v83obus[temp_w*2 +:temp_w];
assign v83ibus[data_w*2 +:data_w] = c1096obus[data_w*0 +:data_w];
assign c1096ibus[temp_w*1 +:temp_w] = v490obus[temp_w*5 +:temp_w];
assign v490ibus[data_w*5 +:data_w] = c1096obus[data_w*1 +:data_w];
assign c1096ibus[temp_w*2 +:temp_w] = v753obus[temp_w*5 +:temp_w];
assign v753ibus[data_w*5 +:data_w] = c1096obus[data_w*2 +:data_w];
assign c1096ibus[temp_w*3 +:temp_w] = v1122obus[temp_w*5 +:temp_w];
assign v1122ibus[data_w*5 +:data_w] = c1096obus[data_w*3 +:data_w];
assign c1096ibus[temp_w*4 +:temp_w] = v1199obus[temp_w*2 +:temp_w];
assign v1199ibus[data_w*2 +:data_w] = c1096obus[data_w*4 +:data_w];
assign c1096ibus[temp_w*5 +:temp_w] = v2248obus[temp_w*1 +:temp_w];
assign v2248ibus[data_w*1 +:data_w] = c1096obus[data_w*5 +:data_w];
assign c1097ibus[temp_w*0 +:temp_w] = v84obus[temp_w*2 +:temp_w];
assign v84ibus[data_w*2 +:data_w] = c1097obus[data_w*0 +:data_w];
assign c1097ibus[temp_w*1 +:temp_w] = v491obus[temp_w*5 +:temp_w];
assign v491ibus[data_w*5 +:data_w] = c1097obus[data_w*1 +:data_w];
assign c1097ibus[temp_w*2 +:temp_w] = v754obus[temp_w*5 +:temp_w];
assign v754ibus[data_w*5 +:data_w] = c1097obus[data_w*2 +:data_w];
assign c1097ibus[temp_w*3 +:temp_w] = v1123obus[temp_w*5 +:temp_w];
assign v1123ibus[data_w*5 +:data_w] = c1097obus[data_w*3 +:data_w];
assign c1097ibus[temp_w*4 +:temp_w] = v1200obus[temp_w*2 +:temp_w];
assign v1200ibus[data_w*2 +:data_w] = c1097obus[data_w*4 +:data_w];
assign c1097ibus[temp_w*5 +:temp_w] = v2249obus[temp_w*1 +:temp_w];
assign v2249ibus[data_w*1 +:data_w] = c1097obus[data_w*5 +:data_w];
assign c1098ibus[temp_w*0 +:temp_w] = v85obus[temp_w*2 +:temp_w];
assign v85ibus[data_w*2 +:data_w] = c1098obus[data_w*0 +:data_w];
assign c1098ibus[temp_w*1 +:temp_w] = v492obus[temp_w*5 +:temp_w];
assign v492ibus[data_w*5 +:data_w] = c1098obus[data_w*1 +:data_w];
assign c1098ibus[temp_w*2 +:temp_w] = v755obus[temp_w*5 +:temp_w];
assign v755ibus[data_w*5 +:data_w] = c1098obus[data_w*2 +:data_w];
assign c1098ibus[temp_w*3 +:temp_w] = v1124obus[temp_w*5 +:temp_w];
assign v1124ibus[data_w*5 +:data_w] = c1098obus[data_w*3 +:data_w];
assign c1098ibus[temp_w*4 +:temp_w] = v1201obus[temp_w*2 +:temp_w];
assign v1201ibus[data_w*2 +:data_w] = c1098obus[data_w*4 +:data_w];
assign c1098ibus[temp_w*5 +:temp_w] = v2250obus[temp_w*1 +:temp_w];
assign v2250ibus[data_w*1 +:data_w] = c1098obus[data_w*5 +:data_w];
assign c1099ibus[temp_w*0 +:temp_w] = v86obus[temp_w*2 +:temp_w];
assign v86ibus[data_w*2 +:data_w] = c1099obus[data_w*0 +:data_w];
assign c1099ibus[temp_w*1 +:temp_w] = v493obus[temp_w*5 +:temp_w];
assign v493ibus[data_w*5 +:data_w] = c1099obus[data_w*1 +:data_w];
assign c1099ibus[temp_w*2 +:temp_w] = v756obus[temp_w*5 +:temp_w];
assign v756ibus[data_w*5 +:data_w] = c1099obus[data_w*2 +:data_w];
assign c1099ibus[temp_w*3 +:temp_w] = v1125obus[temp_w*5 +:temp_w];
assign v1125ibus[data_w*5 +:data_w] = c1099obus[data_w*3 +:data_w];
assign c1099ibus[temp_w*4 +:temp_w] = v1202obus[temp_w*2 +:temp_w];
assign v1202ibus[data_w*2 +:data_w] = c1099obus[data_w*4 +:data_w];
assign c1099ibus[temp_w*5 +:temp_w] = v2251obus[temp_w*1 +:temp_w];
assign v2251ibus[data_w*1 +:data_w] = c1099obus[data_w*5 +:data_w];
assign c1100ibus[temp_w*0 +:temp_w] = v87obus[temp_w*2 +:temp_w];
assign v87ibus[data_w*2 +:data_w] = c1100obus[data_w*0 +:data_w];
assign c1100ibus[temp_w*1 +:temp_w] = v494obus[temp_w*5 +:temp_w];
assign v494ibus[data_w*5 +:data_w] = c1100obus[data_w*1 +:data_w];
assign c1100ibus[temp_w*2 +:temp_w] = v757obus[temp_w*5 +:temp_w];
assign v757ibus[data_w*5 +:data_w] = c1100obus[data_w*2 +:data_w];
assign c1100ibus[temp_w*3 +:temp_w] = v1126obus[temp_w*5 +:temp_w];
assign v1126ibus[data_w*5 +:data_w] = c1100obus[data_w*3 +:data_w];
assign c1100ibus[temp_w*4 +:temp_w] = v1203obus[temp_w*2 +:temp_w];
assign v1203ibus[data_w*2 +:data_w] = c1100obus[data_w*4 +:data_w];
assign c1100ibus[temp_w*5 +:temp_w] = v2252obus[temp_w*1 +:temp_w];
assign v2252ibus[data_w*1 +:data_w] = c1100obus[data_w*5 +:data_w];
assign c1101ibus[temp_w*0 +:temp_w] = v88obus[temp_w*2 +:temp_w];
assign v88ibus[data_w*2 +:data_w] = c1101obus[data_w*0 +:data_w];
assign c1101ibus[temp_w*1 +:temp_w] = v495obus[temp_w*5 +:temp_w];
assign v495ibus[data_w*5 +:data_w] = c1101obus[data_w*1 +:data_w];
assign c1101ibus[temp_w*2 +:temp_w] = v758obus[temp_w*5 +:temp_w];
assign v758ibus[data_w*5 +:data_w] = c1101obus[data_w*2 +:data_w];
assign c1101ibus[temp_w*3 +:temp_w] = v1127obus[temp_w*5 +:temp_w];
assign v1127ibus[data_w*5 +:data_w] = c1101obus[data_w*3 +:data_w];
assign c1101ibus[temp_w*4 +:temp_w] = v1204obus[temp_w*2 +:temp_w];
assign v1204ibus[data_w*2 +:data_w] = c1101obus[data_w*4 +:data_w];
assign c1101ibus[temp_w*5 +:temp_w] = v2253obus[temp_w*1 +:temp_w];
assign v2253ibus[data_w*1 +:data_w] = c1101obus[data_w*5 +:data_w];
assign c1102ibus[temp_w*0 +:temp_w] = v89obus[temp_w*2 +:temp_w];
assign v89ibus[data_w*2 +:data_w] = c1102obus[data_w*0 +:data_w];
assign c1102ibus[temp_w*1 +:temp_w] = v496obus[temp_w*5 +:temp_w];
assign v496ibus[data_w*5 +:data_w] = c1102obus[data_w*1 +:data_w];
assign c1102ibus[temp_w*2 +:temp_w] = v759obus[temp_w*5 +:temp_w];
assign v759ibus[data_w*5 +:data_w] = c1102obus[data_w*2 +:data_w];
assign c1102ibus[temp_w*3 +:temp_w] = v1128obus[temp_w*5 +:temp_w];
assign v1128ibus[data_w*5 +:data_w] = c1102obus[data_w*3 +:data_w];
assign c1102ibus[temp_w*4 +:temp_w] = v1205obus[temp_w*2 +:temp_w];
assign v1205ibus[data_w*2 +:data_w] = c1102obus[data_w*4 +:data_w];
assign c1102ibus[temp_w*5 +:temp_w] = v2254obus[temp_w*1 +:temp_w];
assign v2254ibus[data_w*1 +:data_w] = c1102obus[data_w*5 +:data_w];
assign c1103ibus[temp_w*0 +:temp_w] = v90obus[temp_w*2 +:temp_w];
assign v90ibus[data_w*2 +:data_w] = c1103obus[data_w*0 +:data_w];
assign c1103ibus[temp_w*1 +:temp_w] = v497obus[temp_w*5 +:temp_w];
assign v497ibus[data_w*5 +:data_w] = c1103obus[data_w*1 +:data_w];
assign c1103ibus[temp_w*2 +:temp_w] = v760obus[temp_w*5 +:temp_w];
assign v760ibus[data_w*5 +:data_w] = c1103obus[data_w*2 +:data_w];
assign c1103ibus[temp_w*3 +:temp_w] = v1129obus[temp_w*5 +:temp_w];
assign v1129ibus[data_w*5 +:data_w] = c1103obus[data_w*3 +:data_w];
assign c1103ibus[temp_w*4 +:temp_w] = v1206obus[temp_w*2 +:temp_w];
assign v1206ibus[data_w*2 +:data_w] = c1103obus[data_w*4 +:data_w];
assign c1103ibus[temp_w*5 +:temp_w] = v2255obus[temp_w*1 +:temp_w];
assign v2255ibus[data_w*1 +:data_w] = c1103obus[data_w*5 +:data_w];
assign c1104ibus[temp_w*0 +:temp_w] = v91obus[temp_w*2 +:temp_w];
assign v91ibus[data_w*2 +:data_w] = c1104obus[data_w*0 +:data_w];
assign c1104ibus[temp_w*1 +:temp_w] = v498obus[temp_w*5 +:temp_w];
assign v498ibus[data_w*5 +:data_w] = c1104obus[data_w*1 +:data_w];
assign c1104ibus[temp_w*2 +:temp_w] = v761obus[temp_w*5 +:temp_w];
assign v761ibus[data_w*5 +:data_w] = c1104obus[data_w*2 +:data_w];
assign c1104ibus[temp_w*3 +:temp_w] = v1130obus[temp_w*5 +:temp_w];
assign v1130ibus[data_w*5 +:data_w] = c1104obus[data_w*3 +:data_w];
assign c1104ibus[temp_w*4 +:temp_w] = v1207obus[temp_w*2 +:temp_w];
assign v1207ibus[data_w*2 +:data_w] = c1104obus[data_w*4 +:data_w];
assign c1104ibus[temp_w*5 +:temp_w] = v2256obus[temp_w*1 +:temp_w];
assign v2256ibus[data_w*1 +:data_w] = c1104obus[data_w*5 +:data_w];
assign c1105ibus[temp_w*0 +:temp_w] = v92obus[temp_w*2 +:temp_w];
assign v92ibus[data_w*2 +:data_w] = c1105obus[data_w*0 +:data_w];
assign c1105ibus[temp_w*1 +:temp_w] = v499obus[temp_w*5 +:temp_w];
assign v499ibus[data_w*5 +:data_w] = c1105obus[data_w*1 +:data_w];
assign c1105ibus[temp_w*2 +:temp_w] = v762obus[temp_w*5 +:temp_w];
assign v762ibus[data_w*5 +:data_w] = c1105obus[data_w*2 +:data_w];
assign c1105ibus[temp_w*3 +:temp_w] = v1131obus[temp_w*5 +:temp_w];
assign v1131ibus[data_w*5 +:data_w] = c1105obus[data_w*3 +:data_w];
assign c1105ibus[temp_w*4 +:temp_w] = v1208obus[temp_w*2 +:temp_w];
assign v1208ibus[data_w*2 +:data_w] = c1105obus[data_w*4 +:data_w];
assign c1105ibus[temp_w*5 +:temp_w] = v2257obus[temp_w*1 +:temp_w];
assign v2257ibus[data_w*1 +:data_w] = c1105obus[data_w*5 +:data_w];
assign c1106ibus[temp_w*0 +:temp_w] = v93obus[temp_w*2 +:temp_w];
assign v93ibus[data_w*2 +:data_w] = c1106obus[data_w*0 +:data_w];
assign c1106ibus[temp_w*1 +:temp_w] = v500obus[temp_w*5 +:temp_w];
assign v500ibus[data_w*5 +:data_w] = c1106obus[data_w*1 +:data_w];
assign c1106ibus[temp_w*2 +:temp_w] = v763obus[temp_w*5 +:temp_w];
assign v763ibus[data_w*5 +:data_w] = c1106obus[data_w*2 +:data_w];
assign c1106ibus[temp_w*3 +:temp_w] = v1132obus[temp_w*5 +:temp_w];
assign v1132ibus[data_w*5 +:data_w] = c1106obus[data_w*3 +:data_w];
assign c1106ibus[temp_w*4 +:temp_w] = v1209obus[temp_w*2 +:temp_w];
assign v1209ibus[data_w*2 +:data_w] = c1106obus[data_w*4 +:data_w];
assign c1106ibus[temp_w*5 +:temp_w] = v2258obus[temp_w*1 +:temp_w];
assign v2258ibus[data_w*1 +:data_w] = c1106obus[data_w*5 +:data_w];
assign c1107ibus[temp_w*0 +:temp_w] = v94obus[temp_w*2 +:temp_w];
assign v94ibus[data_w*2 +:data_w] = c1107obus[data_w*0 +:data_w];
assign c1107ibus[temp_w*1 +:temp_w] = v501obus[temp_w*5 +:temp_w];
assign v501ibus[data_w*5 +:data_w] = c1107obus[data_w*1 +:data_w];
assign c1107ibus[temp_w*2 +:temp_w] = v764obus[temp_w*5 +:temp_w];
assign v764ibus[data_w*5 +:data_w] = c1107obus[data_w*2 +:data_w];
assign c1107ibus[temp_w*3 +:temp_w] = v1133obus[temp_w*5 +:temp_w];
assign v1133ibus[data_w*5 +:data_w] = c1107obus[data_w*3 +:data_w];
assign c1107ibus[temp_w*4 +:temp_w] = v1210obus[temp_w*2 +:temp_w];
assign v1210ibus[data_w*2 +:data_w] = c1107obus[data_w*4 +:data_w];
assign c1107ibus[temp_w*5 +:temp_w] = v2259obus[temp_w*1 +:temp_w];
assign v2259ibus[data_w*1 +:data_w] = c1107obus[data_w*5 +:data_w];
assign c1108ibus[temp_w*0 +:temp_w] = v95obus[temp_w*2 +:temp_w];
assign v95ibus[data_w*2 +:data_w] = c1108obus[data_w*0 +:data_w];
assign c1108ibus[temp_w*1 +:temp_w] = v502obus[temp_w*5 +:temp_w];
assign v502ibus[data_w*5 +:data_w] = c1108obus[data_w*1 +:data_w];
assign c1108ibus[temp_w*2 +:temp_w] = v765obus[temp_w*5 +:temp_w];
assign v765ibus[data_w*5 +:data_w] = c1108obus[data_w*2 +:data_w];
assign c1108ibus[temp_w*3 +:temp_w] = v1134obus[temp_w*5 +:temp_w];
assign v1134ibus[data_w*5 +:data_w] = c1108obus[data_w*3 +:data_w];
assign c1108ibus[temp_w*4 +:temp_w] = v1211obus[temp_w*2 +:temp_w];
assign v1211ibus[data_w*2 +:data_w] = c1108obus[data_w*4 +:data_w];
assign c1108ibus[temp_w*5 +:temp_w] = v2260obus[temp_w*1 +:temp_w];
assign v2260ibus[data_w*1 +:data_w] = c1108obus[data_w*5 +:data_w];
assign c1109ibus[temp_w*0 +:temp_w] = v0obus[temp_w*2 +:temp_w];
assign v0ibus[data_w*2 +:data_w] = c1109obus[data_w*0 +:data_w];
assign c1109ibus[temp_w*1 +:temp_w] = v503obus[temp_w*5 +:temp_w];
assign v503ibus[data_w*5 +:data_w] = c1109obus[data_w*1 +:data_w];
assign c1109ibus[temp_w*2 +:temp_w] = v766obus[temp_w*5 +:temp_w];
assign v766ibus[data_w*5 +:data_w] = c1109obus[data_w*2 +:data_w];
assign c1109ibus[temp_w*3 +:temp_w] = v1135obus[temp_w*5 +:temp_w];
assign v1135ibus[data_w*5 +:data_w] = c1109obus[data_w*3 +:data_w];
assign c1109ibus[temp_w*4 +:temp_w] = v1212obus[temp_w*2 +:temp_w];
assign v1212ibus[data_w*2 +:data_w] = c1109obus[data_w*4 +:data_w];
assign c1109ibus[temp_w*5 +:temp_w] = v2261obus[temp_w*1 +:temp_w];
assign v2261ibus[data_w*1 +:data_w] = c1109obus[data_w*5 +:data_w];
assign c1110ibus[temp_w*0 +:temp_w] = v1obus[temp_w*2 +:temp_w];
assign v1ibus[data_w*2 +:data_w] = c1110obus[data_w*0 +:data_w];
assign c1110ibus[temp_w*1 +:temp_w] = v504obus[temp_w*5 +:temp_w];
assign v504ibus[data_w*5 +:data_w] = c1110obus[data_w*1 +:data_w];
assign c1110ibus[temp_w*2 +:temp_w] = v767obus[temp_w*5 +:temp_w];
assign v767ibus[data_w*5 +:data_w] = c1110obus[data_w*2 +:data_w];
assign c1110ibus[temp_w*3 +:temp_w] = v1136obus[temp_w*5 +:temp_w];
assign v1136ibus[data_w*5 +:data_w] = c1110obus[data_w*3 +:data_w];
assign c1110ibus[temp_w*4 +:temp_w] = v1213obus[temp_w*2 +:temp_w];
assign v1213ibus[data_w*2 +:data_w] = c1110obus[data_w*4 +:data_w];
assign c1110ibus[temp_w*5 +:temp_w] = v2262obus[temp_w*1 +:temp_w];
assign v2262ibus[data_w*1 +:data_w] = c1110obus[data_w*5 +:data_w];
assign c1111ibus[temp_w*0 +:temp_w] = v2obus[temp_w*2 +:temp_w];
assign v2ibus[data_w*2 +:data_w] = c1111obus[data_w*0 +:data_w];
assign c1111ibus[temp_w*1 +:temp_w] = v505obus[temp_w*5 +:temp_w];
assign v505ibus[data_w*5 +:data_w] = c1111obus[data_w*1 +:data_w];
assign c1111ibus[temp_w*2 +:temp_w] = v672obus[temp_w*5 +:temp_w];
assign v672ibus[data_w*5 +:data_w] = c1111obus[data_w*2 +:data_w];
assign c1111ibus[temp_w*3 +:temp_w] = v1137obus[temp_w*5 +:temp_w];
assign v1137ibus[data_w*5 +:data_w] = c1111obus[data_w*3 +:data_w];
assign c1111ibus[temp_w*4 +:temp_w] = v1214obus[temp_w*2 +:temp_w];
assign v1214ibus[data_w*2 +:data_w] = c1111obus[data_w*4 +:data_w];
assign c1111ibus[temp_w*5 +:temp_w] = v2263obus[temp_w*1 +:temp_w];
assign v2263ibus[data_w*1 +:data_w] = c1111obus[data_w*5 +:data_w];
assign c1112ibus[temp_w*0 +:temp_w] = v3obus[temp_w*2 +:temp_w];
assign v3ibus[data_w*2 +:data_w] = c1112obus[data_w*0 +:data_w];
assign c1112ibus[temp_w*1 +:temp_w] = v506obus[temp_w*5 +:temp_w];
assign v506ibus[data_w*5 +:data_w] = c1112obus[data_w*1 +:data_w];
assign c1112ibus[temp_w*2 +:temp_w] = v673obus[temp_w*5 +:temp_w];
assign v673ibus[data_w*5 +:data_w] = c1112obus[data_w*2 +:data_w];
assign c1112ibus[temp_w*3 +:temp_w] = v1138obus[temp_w*5 +:temp_w];
assign v1138ibus[data_w*5 +:data_w] = c1112obus[data_w*3 +:data_w];
assign c1112ibus[temp_w*4 +:temp_w] = v1215obus[temp_w*2 +:temp_w];
assign v1215ibus[data_w*2 +:data_w] = c1112obus[data_w*4 +:data_w];
assign c1112ibus[temp_w*5 +:temp_w] = v2264obus[temp_w*1 +:temp_w];
assign v2264ibus[data_w*1 +:data_w] = c1112obus[data_w*5 +:data_w];
assign c1113ibus[temp_w*0 +:temp_w] = v4obus[temp_w*2 +:temp_w];
assign v4ibus[data_w*2 +:data_w] = c1113obus[data_w*0 +:data_w];
assign c1113ibus[temp_w*1 +:temp_w] = v507obus[temp_w*5 +:temp_w];
assign v507ibus[data_w*5 +:data_w] = c1113obus[data_w*1 +:data_w];
assign c1113ibus[temp_w*2 +:temp_w] = v674obus[temp_w*5 +:temp_w];
assign v674ibus[data_w*5 +:data_w] = c1113obus[data_w*2 +:data_w];
assign c1113ibus[temp_w*3 +:temp_w] = v1139obus[temp_w*5 +:temp_w];
assign v1139ibus[data_w*5 +:data_w] = c1113obus[data_w*3 +:data_w];
assign c1113ibus[temp_w*4 +:temp_w] = v1216obus[temp_w*2 +:temp_w];
assign v1216ibus[data_w*2 +:data_w] = c1113obus[data_w*4 +:data_w];
assign c1113ibus[temp_w*5 +:temp_w] = v2265obus[temp_w*1 +:temp_w];
assign v2265ibus[data_w*1 +:data_w] = c1113obus[data_w*5 +:data_w];
assign c1114ibus[temp_w*0 +:temp_w] = v5obus[temp_w*2 +:temp_w];
assign v5ibus[data_w*2 +:data_w] = c1114obus[data_w*0 +:data_w];
assign c1114ibus[temp_w*1 +:temp_w] = v508obus[temp_w*5 +:temp_w];
assign v508ibus[data_w*5 +:data_w] = c1114obus[data_w*1 +:data_w];
assign c1114ibus[temp_w*2 +:temp_w] = v675obus[temp_w*5 +:temp_w];
assign v675ibus[data_w*5 +:data_w] = c1114obus[data_w*2 +:data_w];
assign c1114ibus[temp_w*3 +:temp_w] = v1140obus[temp_w*5 +:temp_w];
assign v1140ibus[data_w*5 +:data_w] = c1114obus[data_w*3 +:data_w];
assign c1114ibus[temp_w*4 +:temp_w] = v1217obus[temp_w*2 +:temp_w];
assign v1217ibus[data_w*2 +:data_w] = c1114obus[data_w*4 +:data_w];
assign c1114ibus[temp_w*5 +:temp_w] = v2266obus[temp_w*1 +:temp_w];
assign v2266ibus[data_w*1 +:data_w] = c1114obus[data_w*5 +:data_w];
assign c1115ibus[temp_w*0 +:temp_w] = v6obus[temp_w*2 +:temp_w];
assign v6ibus[data_w*2 +:data_w] = c1115obus[data_w*0 +:data_w];
assign c1115ibus[temp_w*1 +:temp_w] = v509obus[temp_w*5 +:temp_w];
assign v509ibus[data_w*5 +:data_w] = c1115obus[data_w*1 +:data_w];
assign c1115ibus[temp_w*2 +:temp_w] = v676obus[temp_w*5 +:temp_w];
assign v676ibus[data_w*5 +:data_w] = c1115obus[data_w*2 +:data_w];
assign c1115ibus[temp_w*3 +:temp_w] = v1141obus[temp_w*5 +:temp_w];
assign v1141ibus[data_w*5 +:data_w] = c1115obus[data_w*3 +:data_w];
assign c1115ibus[temp_w*4 +:temp_w] = v1218obus[temp_w*2 +:temp_w];
assign v1218ibus[data_w*2 +:data_w] = c1115obus[data_w*4 +:data_w];
assign c1115ibus[temp_w*5 +:temp_w] = v2267obus[temp_w*1 +:temp_w];
assign v2267ibus[data_w*1 +:data_w] = c1115obus[data_w*5 +:data_w];
assign c1116ibus[temp_w*0 +:temp_w] = v7obus[temp_w*2 +:temp_w];
assign v7ibus[data_w*2 +:data_w] = c1116obus[data_w*0 +:data_w];
assign c1116ibus[temp_w*1 +:temp_w] = v510obus[temp_w*5 +:temp_w];
assign v510ibus[data_w*5 +:data_w] = c1116obus[data_w*1 +:data_w];
assign c1116ibus[temp_w*2 +:temp_w] = v677obus[temp_w*5 +:temp_w];
assign v677ibus[data_w*5 +:data_w] = c1116obus[data_w*2 +:data_w];
assign c1116ibus[temp_w*3 +:temp_w] = v1142obus[temp_w*5 +:temp_w];
assign v1142ibus[data_w*5 +:data_w] = c1116obus[data_w*3 +:data_w];
assign c1116ibus[temp_w*4 +:temp_w] = v1219obus[temp_w*2 +:temp_w];
assign v1219ibus[data_w*2 +:data_w] = c1116obus[data_w*4 +:data_w];
assign c1116ibus[temp_w*5 +:temp_w] = v2268obus[temp_w*1 +:temp_w];
assign v2268ibus[data_w*1 +:data_w] = c1116obus[data_w*5 +:data_w];
assign c1117ibus[temp_w*0 +:temp_w] = v8obus[temp_w*2 +:temp_w];
assign v8ibus[data_w*2 +:data_w] = c1117obus[data_w*0 +:data_w];
assign c1117ibus[temp_w*1 +:temp_w] = v511obus[temp_w*5 +:temp_w];
assign v511ibus[data_w*5 +:data_w] = c1117obus[data_w*1 +:data_w];
assign c1117ibus[temp_w*2 +:temp_w] = v678obus[temp_w*5 +:temp_w];
assign v678ibus[data_w*5 +:data_w] = c1117obus[data_w*2 +:data_w];
assign c1117ibus[temp_w*3 +:temp_w] = v1143obus[temp_w*5 +:temp_w];
assign v1143ibus[data_w*5 +:data_w] = c1117obus[data_w*3 +:data_w];
assign c1117ibus[temp_w*4 +:temp_w] = v1220obus[temp_w*2 +:temp_w];
assign v1220ibus[data_w*2 +:data_w] = c1117obus[data_w*4 +:data_w];
assign c1117ibus[temp_w*5 +:temp_w] = v2269obus[temp_w*1 +:temp_w];
assign v2269ibus[data_w*1 +:data_w] = c1117obus[data_w*5 +:data_w];
assign c1118ibus[temp_w*0 +:temp_w] = v9obus[temp_w*2 +:temp_w];
assign v9ibus[data_w*2 +:data_w] = c1118obus[data_w*0 +:data_w];
assign c1118ibus[temp_w*1 +:temp_w] = v512obus[temp_w*5 +:temp_w];
assign v512ibus[data_w*5 +:data_w] = c1118obus[data_w*1 +:data_w];
assign c1118ibus[temp_w*2 +:temp_w] = v679obus[temp_w*5 +:temp_w];
assign v679ibus[data_w*5 +:data_w] = c1118obus[data_w*2 +:data_w];
assign c1118ibus[temp_w*3 +:temp_w] = v1144obus[temp_w*5 +:temp_w];
assign v1144ibus[data_w*5 +:data_w] = c1118obus[data_w*3 +:data_w];
assign c1118ibus[temp_w*4 +:temp_w] = v1221obus[temp_w*2 +:temp_w];
assign v1221ibus[data_w*2 +:data_w] = c1118obus[data_w*4 +:data_w];
assign c1118ibus[temp_w*5 +:temp_w] = v2270obus[temp_w*1 +:temp_w];
assign v2270ibus[data_w*1 +:data_w] = c1118obus[data_w*5 +:data_w];
assign c1119ibus[temp_w*0 +:temp_w] = v10obus[temp_w*2 +:temp_w];
assign v10ibus[data_w*2 +:data_w] = c1119obus[data_w*0 +:data_w];
assign c1119ibus[temp_w*1 +:temp_w] = v513obus[temp_w*5 +:temp_w];
assign v513ibus[data_w*5 +:data_w] = c1119obus[data_w*1 +:data_w];
assign c1119ibus[temp_w*2 +:temp_w] = v680obus[temp_w*5 +:temp_w];
assign v680ibus[data_w*5 +:data_w] = c1119obus[data_w*2 +:data_w];
assign c1119ibus[temp_w*3 +:temp_w] = v1145obus[temp_w*5 +:temp_w];
assign v1145ibus[data_w*5 +:data_w] = c1119obus[data_w*3 +:data_w];
assign c1119ibus[temp_w*4 +:temp_w] = v1222obus[temp_w*2 +:temp_w];
assign v1222ibus[data_w*2 +:data_w] = c1119obus[data_w*4 +:data_w];
assign c1119ibus[temp_w*5 +:temp_w] = v2271obus[temp_w*1 +:temp_w];
assign v2271ibus[data_w*1 +:data_w] = c1119obus[data_w*5 +:data_w];
assign c1120ibus[temp_w*0 +:temp_w] = v11obus[temp_w*2 +:temp_w];
assign v11ibus[data_w*2 +:data_w] = c1120obus[data_w*0 +:data_w];
assign c1120ibus[temp_w*1 +:temp_w] = v514obus[temp_w*5 +:temp_w];
assign v514ibus[data_w*5 +:data_w] = c1120obus[data_w*1 +:data_w];
assign c1120ibus[temp_w*2 +:temp_w] = v681obus[temp_w*5 +:temp_w];
assign v681ibus[data_w*5 +:data_w] = c1120obus[data_w*2 +:data_w];
assign c1120ibus[temp_w*3 +:temp_w] = v1146obus[temp_w*5 +:temp_w];
assign v1146ibus[data_w*5 +:data_w] = c1120obus[data_w*3 +:data_w];
assign c1120ibus[temp_w*4 +:temp_w] = v1223obus[temp_w*2 +:temp_w];
assign v1223ibus[data_w*2 +:data_w] = c1120obus[data_w*4 +:data_w];
assign c1120ibus[temp_w*5 +:temp_w] = v2272obus[temp_w*1 +:temp_w];
assign v2272ibus[data_w*1 +:data_w] = c1120obus[data_w*5 +:data_w];
assign c1121ibus[temp_w*0 +:temp_w] = v12obus[temp_w*2 +:temp_w];
assign v12ibus[data_w*2 +:data_w] = c1121obus[data_w*0 +:data_w];
assign c1121ibus[temp_w*1 +:temp_w] = v515obus[temp_w*5 +:temp_w];
assign v515ibus[data_w*5 +:data_w] = c1121obus[data_w*1 +:data_w];
assign c1121ibus[temp_w*2 +:temp_w] = v682obus[temp_w*5 +:temp_w];
assign v682ibus[data_w*5 +:data_w] = c1121obus[data_w*2 +:data_w];
assign c1121ibus[temp_w*3 +:temp_w] = v1147obus[temp_w*5 +:temp_w];
assign v1147ibus[data_w*5 +:data_w] = c1121obus[data_w*3 +:data_w];
assign c1121ibus[temp_w*4 +:temp_w] = v1224obus[temp_w*2 +:temp_w];
assign v1224ibus[data_w*2 +:data_w] = c1121obus[data_w*4 +:data_w];
assign c1121ibus[temp_w*5 +:temp_w] = v2273obus[temp_w*1 +:temp_w];
assign v2273ibus[data_w*1 +:data_w] = c1121obus[data_w*5 +:data_w];
assign c1122ibus[temp_w*0 +:temp_w] = v13obus[temp_w*2 +:temp_w];
assign v13ibus[data_w*2 +:data_w] = c1122obus[data_w*0 +:data_w];
assign c1122ibus[temp_w*1 +:temp_w] = v516obus[temp_w*5 +:temp_w];
assign v516ibus[data_w*5 +:data_w] = c1122obus[data_w*1 +:data_w];
assign c1122ibus[temp_w*2 +:temp_w] = v683obus[temp_w*5 +:temp_w];
assign v683ibus[data_w*5 +:data_w] = c1122obus[data_w*2 +:data_w];
assign c1122ibus[temp_w*3 +:temp_w] = v1148obus[temp_w*5 +:temp_w];
assign v1148ibus[data_w*5 +:data_w] = c1122obus[data_w*3 +:data_w];
assign c1122ibus[temp_w*4 +:temp_w] = v1225obus[temp_w*2 +:temp_w];
assign v1225ibus[data_w*2 +:data_w] = c1122obus[data_w*4 +:data_w];
assign c1122ibus[temp_w*5 +:temp_w] = v2274obus[temp_w*1 +:temp_w];
assign v2274ibus[data_w*1 +:data_w] = c1122obus[data_w*5 +:data_w];
assign c1123ibus[temp_w*0 +:temp_w] = v14obus[temp_w*2 +:temp_w];
assign v14ibus[data_w*2 +:data_w] = c1123obus[data_w*0 +:data_w];
assign c1123ibus[temp_w*1 +:temp_w] = v517obus[temp_w*5 +:temp_w];
assign v517ibus[data_w*5 +:data_w] = c1123obus[data_w*1 +:data_w];
assign c1123ibus[temp_w*2 +:temp_w] = v684obus[temp_w*5 +:temp_w];
assign v684ibus[data_w*5 +:data_w] = c1123obus[data_w*2 +:data_w];
assign c1123ibus[temp_w*3 +:temp_w] = v1149obus[temp_w*5 +:temp_w];
assign v1149ibus[data_w*5 +:data_w] = c1123obus[data_w*3 +:data_w];
assign c1123ibus[temp_w*4 +:temp_w] = v1226obus[temp_w*2 +:temp_w];
assign v1226ibus[data_w*2 +:data_w] = c1123obus[data_w*4 +:data_w];
assign c1123ibus[temp_w*5 +:temp_w] = v2275obus[temp_w*1 +:temp_w];
assign v2275ibus[data_w*1 +:data_w] = c1123obus[data_w*5 +:data_w];
assign c1124ibus[temp_w*0 +:temp_w] = v15obus[temp_w*2 +:temp_w];
assign v15ibus[data_w*2 +:data_w] = c1124obus[data_w*0 +:data_w];
assign c1124ibus[temp_w*1 +:temp_w] = v518obus[temp_w*5 +:temp_w];
assign v518ibus[data_w*5 +:data_w] = c1124obus[data_w*1 +:data_w];
assign c1124ibus[temp_w*2 +:temp_w] = v685obus[temp_w*5 +:temp_w];
assign v685ibus[data_w*5 +:data_w] = c1124obus[data_w*2 +:data_w];
assign c1124ibus[temp_w*3 +:temp_w] = v1150obus[temp_w*5 +:temp_w];
assign v1150ibus[data_w*5 +:data_w] = c1124obus[data_w*3 +:data_w];
assign c1124ibus[temp_w*4 +:temp_w] = v1227obus[temp_w*2 +:temp_w];
assign v1227ibus[data_w*2 +:data_w] = c1124obus[data_w*4 +:data_w];
assign c1124ibus[temp_w*5 +:temp_w] = v2276obus[temp_w*1 +:temp_w];
assign v2276ibus[data_w*1 +:data_w] = c1124obus[data_w*5 +:data_w];
assign c1125ibus[temp_w*0 +:temp_w] = v16obus[temp_w*2 +:temp_w];
assign v16ibus[data_w*2 +:data_w] = c1125obus[data_w*0 +:data_w];
assign c1125ibus[temp_w*1 +:temp_w] = v519obus[temp_w*5 +:temp_w];
assign v519ibus[data_w*5 +:data_w] = c1125obus[data_w*1 +:data_w];
assign c1125ibus[temp_w*2 +:temp_w] = v686obus[temp_w*5 +:temp_w];
assign v686ibus[data_w*5 +:data_w] = c1125obus[data_w*2 +:data_w];
assign c1125ibus[temp_w*3 +:temp_w] = v1151obus[temp_w*5 +:temp_w];
assign v1151ibus[data_w*5 +:data_w] = c1125obus[data_w*3 +:data_w];
assign c1125ibus[temp_w*4 +:temp_w] = v1228obus[temp_w*2 +:temp_w];
assign v1228ibus[data_w*2 +:data_w] = c1125obus[data_w*4 +:data_w];
assign c1125ibus[temp_w*5 +:temp_w] = v2277obus[temp_w*1 +:temp_w];
assign v2277ibus[data_w*1 +:data_w] = c1125obus[data_w*5 +:data_w];
assign c1126ibus[temp_w*0 +:temp_w] = v17obus[temp_w*2 +:temp_w];
assign v17ibus[data_w*2 +:data_w] = c1126obus[data_w*0 +:data_w];
assign c1126ibus[temp_w*1 +:temp_w] = v520obus[temp_w*5 +:temp_w];
assign v520ibus[data_w*5 +:data_w] = c1126obus[data_w*1 +:data_w];
assign c1126ibus[temp_w*2 +:temp_w] = v687obus[temp_w*5 +:temp_w];
assign v687ibus[data_w*5 +:data_w] = c1126obus[data_w*2 +:data_w];
assign c1126ibus[temp_w*3 +:temp_w] = v1056obus[temp_w*5 +:temp_w];
assign v1056ibus[data_w*5 +:data_w] = c1126obus[data_w*3 +:data_w];
assign c1126ibus[temp_w*4 +:temp_w] = v1229obus[temp_w*2 +:temp_w];
assign v1229ibus[data_w*2 +:data_w] = c1126obus[data_w*4 +:data_w];
assign c1126ibus[temp_w*5 +:temp_w] = v2278obus[temp_w*1 +:temp_w];
assign v2278ibus[data_w*1 +:data_w] = c1126obus[data_w*5 +:data_w];
assign c1127ibus[temp_w*0 +:temp_w] = v18obus[temp_w*2 +:temp_w];
assign v18ibus[data_w*2 +:data_w] = c1127obus[data_w*0 +:data_w];
assign c1127ibus[temp_w*1 +:temp_w] = v521obus[temp_w*5 +:temp_w];
assign v521ibus[data_w*5 +:data_w] = c1127obus[data_w*1 +:data_w];
assign c1127ibus[temp_w*2 +:temp_w] = v688obus[temp_w*5 +:temp_w];
assign v688ibus[data_w*5 +:data_w] = c1127obus[data_w*2 +:data_w];
assign c1127ibus[temp_w*3 +:temp_w] = v1057obus[temp_w*5 +:temp_w];
assign v1057ibus[data_w*5 +:data_w] = c1127obus[data_w*3 +:data_w];
assign c1127ibus[temp_w*4 +:temp_w] = v1230obus[temp_w*2 +:temp_w];
assign v1230ibus[data_w*2 +:data_w] = c1127obus[data_w*4 +:data_w];
assign c1127ibus[temp_w*5 +:temp_w] = v2279obus[temp_w*1 +:temp_w];
assign v2279ibus[data_w*1 +:data_w] = c1127obus[data_w*5 +:data_w];
assign c1128ibus[temp_w*0 +:temp_w] = v19obus[temp_w*2 +:temp_w];
assign v19ibus[data_w*2 +:data_w] = c1128obus[data_w*0 +:data_w];
assign c1128ibus[temp_w*1 +:temp_w] = v522obus[temp_w*5 +:temp_w];
assign v522ibus[data_w*5 +:data_w] = c1128obus[data_w*1 +:data_w];
assign c1128ibus[temp_w*2 +:temp_w] = v689obus[temp_w*5 +:temp_w];
assign v689ibus[data_w*5 +:data_w] = c1128obus[data_w*2 +:data_w];
assign c1128ibus[temp_w*3 +:temp_w] = v1058obus[temp_w*5 +:temp_w];
assign v1058ibus[data_w*5 +:data_w] = c1128obus[data_w*3 +:data_w];
assign c1128ibus[temp_w*4 +:temp_w] = v1231obus[temp_w*2 +:temp_w];
assign v1231ibus[data_w*2 +:data_w] = c1128obus[data_w*4 +:data_w];
assign c1128ibus[temp_w*5 +:temp_w] = v2280obus[temp_w*1 +:temp_w];
assign v2280ibus[data_w*1 +:data_w] = c1128obus[data_w*5 +:data_w];
assign c1129ibus[temp_w*0 +:temp_w] = v20obus[temp_w*2 +:temp_w];
assign v20ibus[data_w*2 +:data_w] = c1129obus[data_w*0 +:data_w];
assign c1129ibus[temp_w*1 +:temp_w] = v523obus[temp_w*5 +:temp_w];
assign v523ibus[data_w*5 +:data_w] = c1129obus[data_w*1 +:data_w];
assign c1129ibus[temp_w*2 +:temp_w] = v690obus[temp_w*5 +:temp_w];
assign v690ibus[data_w*5 +:data_w] = c1129obus[data_w*2 +:data_w];
assign c1129ibus[temp_w*3 +:temp_w] = v1059obus[temp_w*5 +:temp_w];
assign v1059ibus[data_w*5 +:data_w] = c1129obus[data_w*3 +:data_w];
assign c1129ibus[temp_w*4 +:temp_w] = v1232obus[temp_w*2 +:temp_w];
assign v1232ibus[data_w*2 +:data_w] = c1129obus[data_w*4 +:data_w];
assign c1129ibus[temp_w*5 +:temp_w] = v2281obus[temp_w*1 +:temp_w];
assign v2281ibus[data_w*1 +:data_w] = c1129obus[data_w*5 +:data_w];
assign c1130ibus[temp_w*0 +:temp_w] = v21obus[temp_w*2 +:temp_w];
assign v21ibus[data_w*2 +:data_w] = c1130obus[data_w*0 +:data_w];
assign c1130ibus[temp_w*1 +:temp_w] = v524obus[temp_w*5 +:temp_w];
assign v524ibus[data_w*5 +:data_w] = c1130obus[data_w*1 +:data_w];
assign c1130ibus[temp_w*2 +:temp_w] = v691obus[temp_w*5 +:temp_w];
assign v691ibus[data_w*5 +:data_w] = c1130obus[data_w*2 +:data_w];
assign c1130ibus[temp_w*3 +:temp_w] = v1060obus[temp_w*5 +:temp_w];
assign v1060ibus[data_w*5 +:data_w] = c1130obus[data_w*3 +:data_w];
assign c1130ibus[temp_w*4 +:temp_w] = v1233obus[temp_w*2 +:temp_w];
assign v1233ibus[data_w*2 +:data_w] = c1130obus[data_w*4 +:data_w];
assign c1130ibus[temp_w*5 +:temp_w] = v2282obus[temp_w*1 +:temp_w];
assign v2282ibus[data_w*1 +:data_w] = c1130obus[data_w*5 +:data_w];
assign c1131ibus[temp_w*0 +:temp_w] = v22obus[temp_w*2 +:temp_w];
assign v22ibus[data_w*2 +:data_w] = c1131obus[data_w*0 +:data_w];
assign c1131ibus[temp_w*1 +:temp_w] = v525obus[temp_w*5 +:temp_w];
assign v525ibus[data_w*5 +:data_w] = c1131obus[data_w*1 +:data_w];
assign c1131ibus[temp_w*2 +:temp_w] = v692obus[temp_w*5 +:temp_w];
assign v692ibus[data_w*5 +:data_w] = c1131obus[data_w*2 +:data_w];
assign c1131ibus[temp_w*3 +:temp_w] = v1061obus[temp_w*5 +:temp_w];
assign v1061ibus[data_w*5 +:data_w] = c1131obus[data_w*3 +:data_w];
assign c1131ibus[temp_w*4 +:temp_w] = v1234obus[temp_w*2 +:temp_w];
assign v1234ibus[data_w*2 +:data_w] = c1131obus[data_w*4 +:data_w];
assign c1131ibus[temp_w*5 +:temp_w] = v2283obus[temp_w*1 +:temp_w];
assign v2283ibus[data_w*1 +:data_w] = c1131obus[data_w*5 +:data_w];
assign c1132ibus[temp_w*0 +:temp_w] = v23obus[temp_w*2 +:temp_w];
assign v23ibus[data_w*2 +:data_w] = c1132obus[data_w*0 +:data_w];
assign c1132ibus[temp_w*1 +:temp_w] = v526obus[temp_w*5 +:temp_w];
assign v526ibus[data_w*5 +:data_w] = c1132obus[data_w*1 +:data_w];
assign c1132ibus[temp_w*2 +:temp_w] = v693obus[temp_w*5 +:temp_w];
assign v693ibus[data_w*5 +:data_w] = c1132obus[data_w*2 +:data_w];
assign c1132ibus[temp_w*3 +:temp_w] = v1062obus[temp_w*5 +:temp_w];
assign v1062ibus[data_w*5 +:data_w] = c1132obus[data_w*3 +:data_w];
assign c1132ibus[temp_w*4 +:temp_w] = v1235obus[temp_w*2 +:temp_w];
assign v1235ibus[data_w*2 +:data_w] = c1132obus[data_w*4 +:data_w];
assign c1132ibus[temp_w*5 +:temp_w] = v2284obus[temp_w*1 +:temp_w];
assign v2284ibus[data_w*1 +:data_w] = c1132obus[data_w*5 +:data_w];
assign c1133ibus[temp_w*0 +:temp_w] = v24obus[temp_w*2 +:temp_w];
assign v24ibus[data_w*2 +:data_w] = c1133obus[data_w*0 +:data_w];
assign c1133ibus[temp_w*1 +:temp_w] = v527obus[temp_w*5 +:temp_w];
assign v527ibus[data_w*5 +:data_w] = c1133obus[data_w*1 +:data_w];
assign c1133ibus[temp_w*2 +:temp_w] = v694obus[temp_w*5 +:temp_w];
assign v694ibus[data_w*5 +:data_w] = c1133obus[data_w*2 +:data_w];
assign c1133ibus[temp_w*3 +:temp_w] = v1063obus[temp_w*5 +:temp_w];
assign v1063ibus[data_w*5 +:data_w] = c1133obus[data_w*3 +:data_w];
assign c1133ibus[temp_w*4 +:temp_w] = v1236obus[temp_w*2 +:temp_w];
assign v1236ibus[data_w*2 +:data_w] = c1133obus[data_w*4 +:data_w];
assign c1133ibus[temp_w*5 +:temp_w] = v2285obus[temp_w*1 +:temp_w];
assign v2285ibus[data_w*1 +:data_w] = c1133obus[data_w*5 +:data_w];
assign c1134ibus[temp_w*0 +:temp_w] = v25obus[temp_w*2 +:temp_w];
assign v25ibus[data_w*2 +:data_w] = c1134obus[data_w*0 +:data_w];
assign c1134ibus[temp_w*1 +:temp_w] = v528obus[temp_w*5 +:temp_w];
assign v528ibus[data_w*5 +:data_w] = c1134obus[data_w*1 +:data_w];
assign c1134ibus[temp_w*2 +:temp_w] = v695obus[temp_w*5 +:temp_w];
assign v695ibus[data_w*5 +:data_w] = c1134obus[data_w*2 +:data_w];
assign c1134ibus[temp_w*3 +:temp_w] = v1064obus[temp_w*5 +:temp_w];
assign v1064ibus[data_w*5 +:data_w] = c1134obus[data_w*3 +:data_w];
assign c1134ibus[temp_w*4 +:temp_w] = v1237obus[temp_w*2 +:temp_w];
assign v1237ibus[data_w*2 +:data_w] = c1134obus[data_w*4 +:data_w];
assign c1134ibus[temp_w*5 +:temp_w] = v2286obus[temp_w*1 +:temp_w];
assign v2286ibus[data_w*1 +:data_w] = c1134obus[data_w*5 +:data_w];
assign c1135ibus[temp_w*0 +:temp_w] = v26obus[temp_w*2 +:temp_w];
assign v26ibus[data_w*2 +:data_w] = c1135obus[data_w*0 +:data_w];
assign c1135ibus[temp_w*1 +:temp_w] = v529obus[temp_w*5 +:temp_w];
assign v529ibus[data_w*5 +:data_w] = c1135obus[data_w*1 +:data_w];
assign c1135ibus[temp_w*2 +:temp_w] = v696obus[temp_w*5 +:temp_w];
assign v696ibus[data_w*5 +:data_w] = c1135obus[data_w*2 +:data_w];
assign c1135ibus[temp_w*3 +:temp_w] = v1065obus[temp_w*5 +:temp_w];
assign v1065ibus[data_w*5 +:data_w] = c1135obus[data_w*3 +:data_w];
assign c1135ibus[temp_w*4 +:temp_w] = v1238obus[temp_w*2 +:temp_w];
assign v1238ibus[data_w*2 +:data_w] = c1135obus[data_w*4 +:data_w];
assign c1135ibus[temp_w*5 +:temp_w] = v2287obus[temp_w*1 +:temp_w];
assign v2287ibus[data_w*1 +:data_w] = c1135obus[data_w*5 +:data_w];
assign c1136ibus[temp_w*0 +:temp_w] = v27obus[temp_w*2 +:temp_w];
assign v27ibus[data_w*2 +:data_w] = c1136obus[data_w*0 +:data_w];
assign c1136ibus[temp_w*1 +:temp_w] = v530obus[temp_w*5 +:temp_w];
assign v530ibus[data_w*5 +:data_w] = c1136obus[data_w*1 +:data_w];
assign c1136ibus[temp_w*2 +:temp_w] = v697obus[temp_w*5 +:temp_w];
assign v697ibus[data_w*5 +:data_w] = c1136obus[data_w*2 +:data_w];
assign c1136ibus[temp_w*3 +:temp_w] = v1066obus[temp_w*5 +:temp_w];
assign v1066ibus[data_w*5 +:data_w] = c1136obus[data_w*3 +:data_w];
assign c1136ibus[temp_w*4 +:temp_w] = v1239obus[temp_w*2 +:temp_w];
assign v1239ibus[data_w*2 +:data_w] = c1136obus[data_w*4 +:data_w];
assign c1136ibus[temp_w*5 +:temp_w] = v2288obus[temp_w*1 +:temp_w];
assign v2288ibus[data_w*1 +:data_w] = c1136obus[data_w*5 +:data_w];
assign c1137ibus[temp_w*0 +:temp_w] = v28obus[temp_w*2 +:temp_w];
assign v28ibus[data_w*2 +:data_w] = c1137obus[data_w*0 +:data_w];
assign c1137ibus[temp_w*1 +:temp_w] = v531obus[temp_w*5 +:temp_w];
assign v531ibus[data_w*5 +:data_w] = c1137obus[data_w*1 +:data_w];
assign c1137ibus[temp_w*2 +:temp_w] = v698obus[temp_w*5 +:temp_w];
assign v698ibus[data_w*5 +:data_w] = c1137obus[data_w*2 +:data_w];
assign c1137ibus[temp_w*3 +:temp_w] = v1067obus[temp_w*5 +:temp_w];
assign v1067ibus[data_w*5 +:data_w] = c1137obus[data_w*3 +:data_w];
assign c1137ibus[temp_w*4 +:temp_w] = v1240obus[temp_w*2 +:temp_w];
assign v1240ibus[data_w*2 +:data_w] = c1137obus[data_w*4 +:data_w];
assign c1137ibus[temp_w*5 +:temp_w] = v2289obus[temp_w*1 +:temp_w];
assign v2289ibus[data_w*1 +:data_w] = c1137obus[data_w*5 +:data_w];
assign c1138ibus[temp_w*0 +:temp_w] = v29obus[temp_w*2 +:temp_w];
assign v29ibus[data_w*2 +:data_w] = c1138obus[data_w*0 +:data_w];
assign c1138ibus[temp_w*1 +:temp_w] = v532obus[temp_w*5 +:temp_w];
assign v532ibus[data_w*5 +:data_w] = c1138obus[data_w*1 +:data_w];
assign c1138ibus[temp_w*2 +:temp_w] = v699obus[temp_w*5 +:temp_w];
assign v699ibus[data_w*5 +:data_w] = c1138obus[data_w*2 +:data_w];
assign c1138ibus[temp_w*3 +:temp_w] = v1068obus[temp_w*5 +:temp_w];
assign v1068ibus[data_w*5 +:data_w] = c1138obus[data_w*3 +:data_w];
assign c1138ibus[temp_w*4 +:temp_w] = v1241obus[temp_w*2 +:temp_w];
assign v1241ibus[data_w*2 +:data_w] = c1138obus[data_w*4 +:data_w];
assign c1138ibus[temp_w*5 +:temp_w] = v2290obus[temp_w*1 +:temp_w];
assign v2290ibus[data_w*1 +:data_w] = c1138obus[data_w*5 +:data_w];
assign c1139ibus[temp_w*0 +:temp_w] = v30obus[temp_w*2 +:temp_w];
assign v30ibus[data_w*2 +:data_w] = c1139obus[data_w*0 +:data_w];
assign c1139ibus[temp_w*1 +:temp_w] = v533obus[temp_w*5 +:temp_w];
assign v533ibus[data_w*5 +:data_w] = c1139obus[data_w*1 +:data_w];
assign c1139ibus[temp_w*2 +:temp_w] = v700obus[temp_w*5 +:temp_w];
assign v700ibus[data_w*5 +:data_w] = c1139obus[data_w*2 +:data_w];
assign c1139ibus[temp_w*3 +:temp_w] = v1069obus[temp_w*5 +:temp_w];
assign v1069ibus[data_w*5 +:data_w] = c1139obus[data_w*3 +:data_w];
assign c1139ibus[temp_w*4 +:temp_w] = v1242obus[temp_w*2 +:temp_w];
assign v1242ibus[data_w*2 +:data_w] = c1139obus[data_w*4 +:data_w];
assign c1139ibus[temp_w*5 +:temp_w] = v2291obus[temp_w*1 +:temp_w];
assign v2291ibus[data_w*1 +:data_w] = c1139obus[data_w*5 +:data_w];
assign c1140ibus[temp_w*0 +:temp_w] = v31obus[temp_w*2 +:temp_w];
assign v31ibus[data_w*2 +:data_w] = c1140obus[data_w*0 +:data_w];
assign c1140ibus[temp_w*1 +:temp_w] = v534obus[temp_w*5 +:temp_w];
assign v534ibus[data_w*5 +:data_w] = c1140obus[data_w*1 +:data_w];
assign c1140ibus[temp_w*2 +:temp_w] = v701obus[temp_w*5 +:temp_w];
assign v701ibus[data_w*5 +:data_w] = c1140obus[data_w*2 +:data_w];
assign c1140ibus[temp_w*3 +:temp_w] = v1070obus[temp_w*5 +:temp_w];
assign v1070ibus[data_w*5 +:data_w] = c1140obus[data_w*3 +:data_w];
assign c1140ibus[temp_w*4 +:temp_w] = v1243obus[temp_w*2 +:temp_w];
assign v1243ibus[data_w*2 +:data_w] = c1140obus[data_w*4 +:data_w];
assign c1140ibus[temp_w*5 +:temp_w] = v2292obus[temp_w*1 +:temp_w];
assign v2292ibus[data_w*1 +:data_w] = c1140obus[data_w*5 +:data_w];
assign c1141ibus[temp_w*0 +:temp_w] = v32obus[temp_w*2 +:temp_w];
assign v32ibus[data_w*2 +:data_w] = c1141obus[data_w*0 +:data_w];
assign c1141ibus[temp_w*1 +:temp_w] = v535obus[temp_w*5 +:temp_w];
assign v535ibus[data_w*5 +:data_w] = c1141obus[data_w*1 +:data_w];
assign c1141ibus[temp_w*2 +:temp_w] = v702obus[temp_w*5 +:temp_w];
assign v702ibus[data_w*5 +:data_w] = c1141obus[data_w*2 +:data_w];
assign c1141ibus[temp_w*3 +:temp_w] = v1071obus[temp_w*5 +:temp_w];
assign v1071ibus[data_w*5 +:data_w] = c1141obus[data_w*3 +:data_w];
assign c1141ibus[temp_w*4 +:temp_w] = v1244obus[temp_w*2 +:temp_w];
assign v1244ibus[data_w*2 +:data_w] = c1141obus[data_w*4 +:data_w];
assign c1141ibus[temp_w*5 +:temp_w] = v2293obus[temp_w*1 +:temp_w];
assign v2293ibus[data_w*1 +:data_w] = c1141obus[data_w*5 +:data_w];
assign c1142ibus[temp_w*0 +:temp_w] = v33obus[temp_w*2 +:temp_w];
assign v33ibus[data_w*2 +:data_w] = c1142obus[data_w*0 +:data_w];
assign c1142ibus[temp_w*1 +:temp_w] = v536obus[temp_w*5 +:temp_w];
assign v536ibus[data_w*5 +:data_w] = c1142obus[data_w*1 +:data_w];
assign c1142ibus[temp_w*2 +:temp_w] = v703obus[temp_w*5 +:temp_w];
assign v703ibus[data_w*5 +:data_w] = c1142obus[data_w*2 +:data_w];
assign c1142ibus[temp_w*3 +:temp_w] = v1072obus[temp_w*5 +:temp_w];
assign v1072ibus[data_w*5 +:data_w] = c1142obus[data_w*3 +:data_w];
assign c1142ibus[temp_w*4 +:temp_w] = v1245obus[temp_w*2 +:temp_w];
assign v1245ibus[data_w*2 +:data_w] = c1142obus[data_w*4 +:data_w];
assign c1142ibus[temp_w*5 +:temp_w] = v2294obus[temp_w*1 +:temp_w];
assign v2294ibus[data_w*1 +:data_w] = c1142obus[data_w*5 +:data_w];
assign c1143ibus[temp_w*0 +:temp_w] = v34obus[temp_w*2 +:temp_w];
assign v34ibus[data_w*2 +:data_w] = c1143obus[data_w*0 +:data_w];
assign c1143ibus[temp_w*1 +:temp_w] = v537obus[temp_w*5 +:temp_w];
assign v537ibus[data_w*5 +:data_w] = c1143obus[data_w*1 +:data_w];
assign c1143ibus[temp_w*2 +:temp_w] = v704obus[temp_w*5 +:temp_w];
assign v704ibus[data_w*5 +:data_w] = c1143obus[data_w*2 +:data_w];
assign c1143ibus[temp_w*3 +:temp_w] = v1073obus[temp_w*5 +:temp_w];
assign v1073ibus[data_w*5 +:data_w] = c1143obus[data_w*3 +:data_w];
assign c1143ibus[temp_w*4 +:temp_w] = v1246obus[temp_w*2 +:temp_w];
assign v1246ibus[data_w*2 +:data_w] = c1143obus[data_w*4 +:data_w];
assign c1143ibus[temp_w*5 +:temp_w] = v2295obus[temp_w*1 +:temp_w];
assign v2295ibus[data_w*1 +:data_w] = c1143obus[data_w*5 +:data_w];
assign c1144ibus[temp_w*0 +:temp_w] = v35obus[temp_w*2 +:temp_w];
assign v35ibus[data_w*2 +:data_w] = c1144obus[data_w*0 +:data_w];
assign c1144ibus[temp_w*1 +:temp_w] = v538obus[temp_w*5 +:temp_w];
assign v538ibus[data_w*5 +:data_w] = c1144obus[data_w*1 +:data_w];
assign c1144ibus[temp_w*2 +:temp_w] = v705obus[temp_w*5 +:temp_w];
assign v705ibus[data_w*5 +:data_w] = c1144obus[data_w*2 +:data_w];
assign c1144ibus[temp_w*3 +:temp_w] = v1074obus[temp_w*5 +:temp_w];
assign v1074ibus[data_w*5 +:data_w] = c1144obus[data_w*3 +:data_w];
assign c1144ibus[temp_w*4 +:temp_w] = v1247obus[temp_w*2 +:temp_w];
assign v1247ibus[data_w*2 +:data_w] = c1144obus[data_w*4 +:data_w];
assign c1144ibus[temp_w*5 +:temp_w] = v2296obus[temp_w*1 +:temp_w];
assign v2296ibus[data_w*1 +:data_w] = c1144obus[data_w*5 +:data_w];
assign c1145ibus[temp_w*0 +:temp_w] = v36obus[temp_w*2 +:temp_w];
assign v36ibus[data_w*2 +:data_w] = c1145obus[data_w*0 +:data_w];
assign c1145ibus[temp_w*1 +:temp_w] = v539obus[temp_w*5 +:temp_w];
assign v539ibus[data_w*5 +:data_w] = c1145obus[data_w*1 +:data_w];
assign c1145ibus[temp_w*2 +:temp_w] = v706obus[temp_w*5 +:temp_w];
assign v706ibus[data_w*5 +:data_w] = c1145obus[data_w*2 +:data_w];
assign c1145ibus[temp_w*3 +:temp_w] = v1075obus[temp_w*5 +:temp_w];
assign v1075ibus[data_w*5 +:data_w] = c1145obus[data_w*3 +:data_w];
assign c1145ibus[temp_w*4 +:temp_w] = v1152obus[temp_w*2 +:temp_w];
assign v1152ibus[data_w*2 +:data_w] = c1145obus[data_w*4 +:data_w];
assign c1145ibus[temp_w*5 +:temp_w] = v2297obus[temp_w*1 +:temp_w];
assign v2297ibus[data_w*1 +:data_w] = c1145obus[data_w*5 +:data_w];
assign c1146ibus[temp_w*0 +:temp_w] = v37obus[temp_w*2 +:temp_w];
assign v37ibus[data_w*2 +:data_w] = c1146obus[data_w*0 +:data_w];
assign c1146ibus[temp_w*1 +:temp_w] = v540obus[temp_w*5 +:temp_w];
assign v540ibus[data_w*5 +:data_w] = c1146obus[data_w*1 +:data_w];
assign c1146ibus[temp_w*2 +:temp_w] = v707obus[temp_w*5 +:temp_w];
assign v707ibus[data_w*5 +:data_w] = c1146obus[data_w*2 +:data_w];
assign c1146ibus[temp_w*3 +:temp_w] = v1076obus[temp_w*5 +:temp_w];
assign v1076ibus[data_w*5 +:data_w] = c1146obus[data_w*3 +:data_w];
assign c1146ibus[temp_w*4 +:temp_w] = v1153obus[temp_w*2 +:temp_w];
assign v1153ibus[data_w*2 +:data_w] = c1146obus[data_w*4 +:data_w];
assign c1146ibus[temp_w*5 +:temp_w] = v2298obus[temp_w*1 +:temp_w];
assign v2298ibus[data_w*1 +:data_w] = c1146obus[data_w*5 +:data_w];
assign c1147ibus[temp_w*0 +:temp_w] = v38obus[temp_w*2 +:temp_w];
assign v38ibus[data_w*2 +:data_w] = c1147obus[data_w*0 +:data_w];
assign c1147ibus[temp_w*1 +:temp_w] = v541obus[temp_w*5 +:temp_w];
assign v541ibus[data_w*5 +:data_w] = c1147obus[data_w*1 +:data_w];
assign c1147ibus[temp_w*2 +:temp_w] = v708obus[temp_w*5 +:temp_w];
assign v708ibus[data_w*5 +:data_w] = c1147obus[data_w*2 +:data_w];
assign c1147ibus[temp_w*3 +:temp_w] = v1077obus[temp_w*5 +:temp_w];
assign v1077ibus[data_w*5 +:data_w] = c1147obus[data_w*3 +:data_w];
assign c1147ibus[temp_w*4 +:temp_w] = v1154obus[temp_w*2 +:temp_w];
assign v1154ibus[data_w*2 +:data_w] = c1147obus[data_w*4 +:data_w];
assign c1147ibus[temp_w*5 +:temp_w] = v2299obus[temp_w*1 +:temp_w];
assign v2299ibus[data_w*1 +:data_w] = c1147obus[data_w*5 +:data_w];
assign c1148ibus[temp_w*0 +:temp_w] = v39obus[temp_w*2 +:temp_w];
assign v39ibus[data_w*2 +:data_w] = c1148obus[data_w*0 +:data_w];
assign c1148ibus[temp_w*1 +:temp_w] = v542obus[temp_w*5 +:temp_w];
assign v542ibus[data_w*5 +:data_w] = c1148obus[data_w*1 +:data_w];
assign c1148ibus[temp_w*2 +:temp_w] = v709obus[temp_w*5 +:temp_w];
assign v709ibus[data_w*5 +:data_w] = c1148obus[data_w*2 +:data_w];
assign c1148ibus[temp_w*3 +:temp_w] = v1078obus[temp_w*5 +:temp_w];
assign v1078ibus[data_w*5 +:data_w] = c1148obus[data_w*3 +:data_w];
assign c1148ibus[temp_w*4 +:temp_w] = v1155obus[temp_w*2 +:temp_w];
assign v1155ibus[data_w*2 +:data_w] = c1148obus[data_w*4 +:data_w];
assign c1148ibus[temp_w*5 +:temp_w] = v2300obus[temp_w*1 +:temp_w];
assign v2300ibus[data_w*1 +:data_w] = c1148obus[data_w*5 +:data_w];
assign c1149ibus[temp_w*0 +:temp_w] = v40obus[temp_w*2 +:temp_w];
assign v40ibus[data_w*2 +:data_w] = c1149obus[data_w*0 +:data_w];
assign c1149ibus[temp_w*1 +:temp_w] = v543obus[temp_w*5 +:temp_w];
assign v543ibus[data_w*5 +:data_w] = c1149obus[data_w*1 +:data_w];
assign c1149ibus[temp_w*2 +:temp_w] = v710obus[temp_w*5 +:temp_w];
assign v710ibus[data_w*5 +:data_w] = c1149obus[data_w*2 +:data_w];
assign c1149ibus[temp_w*3 +:temp_w] = v1079obus[temp_w*5 +:temp_w];
assign v1079ibus[data_w*5 +:data_w] = c1149obus[data_w*3 +:data_w];
assign c1149ibus[temp_w*4 +:temp_w] = v1156obus[temp_w*2 +:temp_w];
assign v1156ibus[data_w*2 +:data_w] = c1149obus[data_w*4 +:data_w];
assign c1149ibus[temp_w*5 +:temp_w] = v2301obus[temp_w*1 +:temp_w];
assign v2301ibus[data_w*1 +:data_w] = c1149obus[data_w*5 +:data_w];
assign c1150ibus[temp_w*0 +:temp_w] = v41obus[temp_w*2 +:temp_w];
assign v41ibus[data_w*2 +:data_w] = c1150obus[data_w*0 +:data_w];
assign c1150ibus[temp_w*1 +:temp_w] = v544obus[temp_w*5 +:temp_w];
assign v544ibus[data_w*5 +:data_w] = c1150obus[data_w*1 +:data_w];
assign c1150ibus[temp_w*2 +:temp_w] = v711obus[temp_w*5 +:temp_w];
assign v711ibus[data_w*5 +:data_w] = c1150obus[data_w*2 +:data_w];
assign c1150ibus[temp_w*3 +:temp_w] = v1080obus[temp_w*5 +:temp_w];
assign v1080ibus[data_w*5 +:data_w] = c1150obus[data_w*3 +:data_w];
assign c1150ibus[temp_w*4 +:temp_w] = v1157obus[temp_w*2 +:temp_w];
assign v1157ibus[data_w*2 +:data_w] = c1150obus[data_w*4 +:data_w];
assign c1150ibus[temp_w*5 +:temp_w] = v2302obus[temp_w*1 +:temp_w];
assign v2302ibus[data_w*1 +:data_w] = c1150obus[data_w*5 +:data_w];
assign c1151ibus[temp_w*0 +:temp_w] = v42obus[temp_w*2 +:temp_w];
assign v42ibus[data_w*2 +:data_w] = c1151obus[data_w*0 +:data_w];
assign c1151ibus[temp_w*1 +:temp_w] = v545obus[temp_w*5 +:temp_w];
assign v545ibus[data_w*5 +:data_w] = c1151obus[data_w*1 +:data_w];
assign c1151ibus[temp_w*2 +:temp_w] = v712obus[temp_w*5 +:temp_w];
assign v712ibus[data_w*5 +:data_w] = c1151obus[data_w*2 +:data_w];
assign c1151ibus[temp_w*3 +:temp_w] = v1081obus[temp_w*5 +:temp_w];
assign v1081ibus[data_w*5 +:data_w] = c1151obus[data_w*3 +:data_w];
assign c1151ibus[temp_w*4 +:temp_w] = v1158obus[temp_w*2 +:temp_w];
assign v1158ibus[data_w*2 +:data_w] = c1151obus[data_w*4 +:data_w];
assign c1151ibus[temp_w*5 +:temp_w] = v2303obus[temp_w*1 +:temp_w];
assign v2303ibus[data_w*1 +:data_w] = c1151obus[data_w*5 +:data_w];

endmodule
