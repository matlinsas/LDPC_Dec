module t;
wire [16*2304-1:0] sig;
reg llr_in;
wire signed [4:0] llr [2303:0];
genvar i;
integer j;

/*
initial begin
    #1000
    for(j=0; j<2304; j=j+1)
        $write("%d ", llr[j]);
end

generate
for(i=0; i<2304; i=i+1) begin :test
    quant Q(
        .snr_idx(4'd10),
        .frac_w(-5'd1),
        .data_in(sig[i*16 +:16]),
        .llr(llr[i])
    );
end
endgenerate 

assign sig = {16'd2224,-16'd4003,-16'd1083,16'd3317,-16'd4628,16'd287,16'd2037,16'd3670,-16'd157,-16'd494,-16'd4171,16'd546,-16'd1630,-16'd1565,16'd665,-16'd326,-16'd1251,-16'd2509,16'd209,-16'd1792,-16'd1604,16'd793,16'd2632,-16'd750,16'd329,-16'd980,16'd25,-16'd2036,-16'd1841,-16'd798,16'd2867,-16'd1579,-16'd961,16'd2886,-16'd2103,16'd1203,-16'd1682,-16'd122,16'd446,16'd1331,-16'd372,-16'd1368,-16'd450,16'd2414,16'd3918,16'd667,16'd2293,-16'd1699,16'd588,16'd2351,16'd176,-16'd786,-16'd2508,16'd3581,16'd434,16'd1600,16'd3423,-16'd335,-16'd1676,-16'd156,-16'd3420,-16'd1992,16'd316,-16'd367,16'd3474,16'd1580,16'd343,16'd893,16'd650,16'd535,-16'd76,-16'd1841,16'd1591,16'd499,-16'd2310,-16'd1477,-16'd597,-16'd1874,16'd431,16'd182,-16'd2123,16'd3775,-16'd4100,-16'd955,16'd1709,16'd3430,-16'd2151,-16'd1249,16'd3661,16'd716,-16'd1949,16'd585,-16'd3239,-16'd3209,16'd1201,-16'd3762,-16'd780,16'd2458,-16'd1890,16'd4737,16'd2380,-16'd3327,16'd2018,-16'd3031,-16'd2320,16'd3933,16'd2075,16'd4159,16'd2567,16'd558,16'd3153,-16'd3484,16'd1058,-16'd891,16'd122,16'd2293,16'd3284,-16'd1006,-16'd1938,-16'd437,16'd1494,-16'd298,-16'd190,16'd1505,-16'd1399,16'd1848,16'd1405,-16'd497,16'd3675,-16'd3758,16'd2994,-16'd58,-16'd2599,16'd626,-16'd2418,16'd4910,16'd1284,-16'd3889,-16'd1540,-16'd18,-16'd959,16'd1050,-16'd3984,16'd2094,-16'd3290,-16'd2254,-16'd1552,16'd5216,-16'd894,16'd2755,-16'd2074,-16'd209,16'd3223,-16'd1082,16'd1614,16'd1677,16'd1024,-16'd1985,-16'd664,16'd1235,-16'd766,-16'd838,16'd3991,16'd1479,16'd703,-16'd1912,16'd1124,-16'd3443,16'd1579,16'd1332,16'd394,16'd3198,-16'd1624,16'd3721,-16'd52,-16'd1049,16'd3354,-16'd3842,-16'd2378,-16'd143,16'd2699,16'd1108,16'd957,-16'd881,-16'd6490,-16'd3310,16'd152,16'd3,16'd2331,16'd1082,16'd1668,16'd832,-16'd726,16'd946,16'd1295,-16'd831,16'd589,16'd1823,-16'd625,-16'd1687,16'd4040,-16'd1641,16'd6107,16'd289,-16'd1667,-16'd1265,-16'd1780,16'd695,-16'd641,-16'd828,-16'd307,16'd1518,16'd1903,-16'd1566,-16'd3195,-16'd2416,-16'd2046,-16'd1400,-16'd2616,-16'd1334,16'd478,16'd1270,16'd103,16'd1267,-16'd1805,-16'd1244,-16'd781,-16'd1654,-16'd734,-16'd325,-16'd2327,16'd3750,16'd2738,16'd2803,16'd1846,-16'd1655,16'd837,16'd243,16'd1021,16'd3296,-16'd1204,16'd2200,16'd1160,16'd1042,-16'd309,-16'd2674,-16'd875,-16'd1841,-16'd736,16'd3653,-16'd3200,-16'd1448,16'd1945,-16'd2538,16'd2429,16'd1390,16'd2148,16'd3362,16'd1848,-16'd3825,16'd160,16'd1737,-16'd5944,-16'd1445,-16'd275,-16'd115,16'd2579,-16'd916,-16'd924,-16'd796,-16'd582,-16'd3892,16'd1649,16'd29,16'd546,-16'd56,-16'd1314,16'd243,16'd3998,16'd895,-16'd32,16'd3018,16'd1583,-16'd473,-16'd1092,-16'd1342,-16'd1144,-16'd3604,-16'd865,-16'd1913,16'd7881,-16'd3147,-16'd454,-16'd1439,-16'd312,16'd595,16'd2607,16'd2988,-16'd1531,16'd278,-16'd1133,-16'd1669,16'd2623,16'd2819,-16'd323,16'd18,-16'd1494,16'd1007,-16'd2047,-16'd3494,16'd2239,16'd884,16'd106,16'd1843,-16'd267,-16'd2193,16'd2616,-16'd4504,16'd260,16'd4662,-16'd2822,16'd13,-16'd1280,16'd3430,-16'd119,16'd953,-16'd775,-16'd447,16'd4180,16'd1773,16'd3548,-16'd101,16'd201,16'd1868,16'd1051,-16'd1481,-16'd1830,-16'd169,16'd766,16'd616,16'd699,16'd3723,16'd3371,16'd2576,-16'd165,16'd1719,-16'd3795,16'd1029,-16'd2127,-16'd2623,-16'd1160,16'd3691,16'd3232,16'd880,16'd4096,16'd1350,-16'd1327,16'd132,-16'd142,-16'd215,16'd2719,16'd387,-16'd3469,16'd3904,16'd1173,16'd3145,16'd844,16'd489,16'd3572,-16'd3288,-16'd1496,16'd993,-16'd3316,16'd759,16'd1174,-16'd420,-16'd673,-16'd2087,-16'd1077,16'd1134,16'd781,-16'd2171,16'd846,-16'd924,-16'd2608,-16'd2678,-16'd2042,16'd1041,-16'd3065,-16'd2093,-16'd298,-16'd4732,-16'd1443,16'd4128,16'd382,16'd1076,16'd2899,-16'd6048,-16'd2338,-16'd4185,16'd3399,-16'd1598,-16'd111,-16'd507,-16'd1211,-16'd152,16'd1865,-16'd426,-16'd383,-16'd2816,16'd1879,16'd5457,-16'd1431,16'd1247,16'd4489,16'd2933,16'd1004,16'd3153,-16'd3862,16'd174,16'd3538,-16'd1850,-16'd2444,-16'd1801,-16'd1822,16'd518,-16'd945,16'd660,-16'd961,16'd1265,-16'd1048,16'd722,16'd984,-16'd2741,16'd1568,16'd599,16'd2429,16'd2166,16'd3793,16'd1214,16'd2451,-16'd1212,16'd2682,16'd3350,-16'd1251,-16'd657,16'd3836,16'd589,-16'd4786,16'd4942,-16'd1278,16'd3817,-16'd643,16'd1156,16'd3647,-16'd109,-16'd4795,-16'd74,16'd265,16'd491,16'd502,16'd521,-16'd319,-16'd1367,-16'd3139,16'd2887,-16'd1689,-16'd2694,16'd1719,-16'd965,16'd2321,16'd2771,-16'd4165,16'd1658,16'd3140,16'd1841,16'd1721,16'd1254,16'd999,16'd2675,16'd434,16'd2906,-16'd1976,16'd2690,-16'd71,16'd3309,-16'd2491,-16'd865,-16'd2048,16'd123,16'd1202,-16'd3249,-16'd2624,16'd4145,16'd1450,16'd799,-16'd3546,-16'd2315,16'd1210,-16'd590,16'd2266,16'd3717,-16'd5189,16'd2208,-16'd650,-16'd1598,16'd2253,-16'd2538,-16'd80,16'd1556,16'd3281,16'd1512,-16'd1587,16'd3821,16'd847,16'd759,16'd1035,-16'd2743,16'd990,16'd3939,16'd2306,-16'd682,-16'd1195,-16'd4090,16'd1717,-16'd1240,-16'd1854,16'd1445,16'd751,16'd59,16'd1674,16'd1429,-16'd1947,-16'd2664,-16'd383,16'd2836,16'd748,-16'd1951,-16'd616,-16'd4819,-16'd928,-16'd3085,-16'd671,-16'd1970,-16'd477,-16'd2973,-16'd477,-16'd180,-16'd353,-16'd2033,-16'd1369,16'd1651,16'd561,-16'd2621,-16'd1007,16'd705,16'd191,16'd4827,-16'd2624,16'd2302,-16'd1574,16'd2453,16'd2907,-16'd87,-16'd317,16'd585,16'd3745,-16'd2196,16'd1582,-16'd1351,16'd563,-16'd1112,-16'd1490,-16'd3779,16'd2959,-16'd2292,16'd1774,-16'd902,16'd1075,16'd925,-16'd2506,-16'd289,-16'd2391,-16'd1496,16'd361,-16'd1428,-16'd2161,-16'd3997,-16'd650,16'd2926,16'd2746,-16'd455,16'd927,-16'd440,-16'd1354,16'd553,-16'd545,16'd1429,16'd1741,-16'd549,-16'd1323,-16'd2410,16'd884,16'd646,16'd1001,16'd3347,16'd1972,-16'd1179,16'd1095,16'd1300,16'd1673,-16'd20,16'd1798,16'd348,-16'd955,16'd2249,-16'd2516,-16'd2677,16'd816,-16'd558,16'd582,16'd234,16'd3997,-16'd2954,-16'd2507,16'd3789,-16'd1122,-16'd1052,16'd213,16'd1128,-16'd1520,16'd139,-16'd3315,16'd621,-16'd1117,-16'd25,-16'd301,16'd1741,16'd3238,16'd2856,-16'd1362,16'd1848,-16'd1108,16'd176,-16'd3471,-16'd489,-16'd971,16'd841,-16'd705,16'd968,16'd2192,16'd1943,16'd409,16'd1023,-16'd1625,-16'd1604,-16'd3112,16'd723,-16'd60,-16'd906,16'd134,-16'd1514,-16'd2885,16'd1559,16'd475,-16'd606,16'd1441,-16'd4104,16'd683,-16'd25,-16'd345,16'd1140,16'd3489,16'd1500,16'd2430,-16'd2676,16'd799,16'd143,-16'd356,-16'd605,16'd1037,16'd1374,16'd1041,16'd1345,16'd538,-16'd841,-16'd697,-16'd114,-16'd2104,-16'd532,16'd514,16'd221,-16'd679,16'd136,-16'd1034,-16'd1008,-16'd96,16'd278,-16'd566,16'd15,-16'd543,-16'd2774,16'd3928,-16'd721,16'd835,16'd622,16'd1151,16'd437,16'd936,16'd783,-16'd264,-16'd2959,-16'd2166,-16'd496,16'd3231,16'd1717,16'd925,16'd230,16'd1058,16'd429,16'd1393,-16'd4177,-16'd1207,16'd842,-16'd864,16'd558,16'd2616,-16'd1676,16'd2558,16'd1168,-16'd493,-16'd428,-16'd4413,16'd1643,16'd3025,16'd1720,-16'd2281,-16'd1015,-16'd1992,-16'd3073,-16'd1390,16'd2289,16'd402,-16'd862,16'd2322,-16'd1373,16'd1927,-16'd1537,16'd468,16'd1531,-16'd1436,16'd2291,16'd2561,16'd1353,-16'd1002,16'd599,16'd2892,-16'd34,-16'd2954,-16'd193,-16'd1989,16'd1505,16'd77,-16'd3165,-16'd443,16'd2761,16'd1562,16'd1133,-16'd3258,-16'd1257,16'd2180,16'd1063,-16'd263,16'd1214,16'd813,-16'd2175,-16'd874,-16'd4417,16'd3229,-16'd2582,-16'd1391,16'd945,-16'd1636,16'd106,-16'd1503,16'd279,-16'd132,16'd2492,-16'd1810,16'd2394,-16'd403,16'd2458,-16'd607,16'd3411,-16'd116,16'd259,-16'd3008,16'd313,-16'd1853,16'd1395,16'd146,-16'd1086,16'd3246,-16'd554,-16'd1611,-16'd255,16'd430,-16'd1534,-16'd2193,-16'd2910,-16'd242,-16'd1744,-16'd689,16'd586,16'd2178,16'd2457,-16'd130,16'd1309,-16'd3738,16'd999,16'd540,-16'd730,16'd1647,-16'd1943,16'd1043,-16'd802,-16'd3741,16'd1461,16'd188,-16'd2570,-16'd417,-16'd26,-16'd301,16'd1710,-16'd1049,16'd2370,16'd1899,-16'd1788,16'd82,-16'd62,-16'd1640,-16'd199,-16'd425,-16'd2816,16'd4753,16'd745,16'd113,16'd2057,-16'd3941,16'd3815,-16'd6337,-16'd1682,-16'd1,-16'd3826,-16'd1524,16'd2787,16'd203,16'd928,16'd215,16'd1515,-16'd469,-16'd2880,16'd1537,-16'd1587,-16'd1755,-16'd3272,-16'd497,16'd4047,16'd175,-16'd2369,-16'd934,-16'd47,16'd1209,-16'd2580,16'd429,16'd6052,-16'd449,16'd18,-16'd784,-16'd2068,16'd1211,16'd983,-16'd468,16'd783,-16'd1010,-16'd1094,16'd485,-16'd3778,16'd3073,16'd1424,-16'd682,-16'd1642,16'd668,16'd4476,16'd680,-16'd2457,16'd3462,-16'd1566,-16'd1797,-16'd530,-16'd722,-16'd659,-16'd1387,-16'd2766,16'd959,16'd644,-16'd970,16'd1815,16'd5258,-16'd245,-16'd2476,16'd596,16'd3081,16'd3260,16'd782,-16'd359,-16'd4157,16'd4110,16'd226,-16'd844,16'd381,16'd2526,-16'd143,16'd731,16'd2529,-16'd2155,-16'd1109,-16'd82,16'd1556,-16'd594,-16'd2609,16'd2506,-16'd1468,-16'd985,16'd2466,16'd1988,16'd479,-16'd29,-16'd3528,-16'd1598,-16'd274,16'd51,16'd551,-16'd113,-16'd385,16'd34,-16'd1951,-16'd302,-16'd1999,16'd898,16'd355,-16'd2687,-16'd1129,16'd2224,-16'd1994,16'd3583,16'd1310,-16'd2695,16'd3314,-16'd4073,16'd1859,16'd987,16'd928,16'd3963,-16'd1686,16'd792,-16'd98,-16'd1244,-16'd3519,16'd2324,16'd961,16'd1092,16'd2208,-16'd509,16'd731,16'd1531,16'd470,16'd2915,-16'd2617,16'd728,-16'd2091,-16'd2548,-16'd1735,16'd1445,-16'd2511,16'd2328,16'd499,-16'd1701,16'd2261,-16'd1179,-16'd779,16'd652,-16'd173,16'd3432,-16'd1116,16'd2957,16'd916,16'd1099,-16'd714,16'd2425,16'd422,16'd271,-16'd1071,16'd1925,-16'd2790,-16'd1622,16'd1358,16'd1199,-16'd444,-16'd1425,-16'd3165,16'd7462,-16'd1574,-16'd433,-16'd1537,16'd405,-16'd298,-16'd3577,-16'd3195,-16'd1195,16'd3132,-16'd930,16'd1169,16'd1393,16'd2460,16'd1692,16'd1270,16'd1160,16'd463,16'd4791,16'd1198,-16'd510,-16'd734,16'd2758,16'd1641,-16'd1117,-16'd410,-16'd1882,-16'd846,16'd337,-16'd1306,-16'd1184,-16'd2166,16'd763,-16'd413,-16'd2981,16'd963,16'd1750,-16'd2804,-16'd1999,-16'd1466,-16'd6045,16'd337,16'd1418,16'd2597,16'd3690,-16'd1652,-16'd2822,-16'd1387,16'd2651,16'd862,-16'd1351,-16'd3204,16'd1739,-16'd534,-16'd2304,16'd776,-16'd895,16'd937,-16'd1742,16'd2284,-16'd1673,16'd237,-16'd1156,16'd1720,-16'd896,16'd2735,-16'd2150,16'd2776,16'd545,16'd754,-16'd2159,16'd645,16'd3655,16'd1928,-16'd810,16'd1471,-16'd1329,-16'd364,16'd2260,16'd92,16'd1776,-16'd812,-16'd1104,16'd2700,-16'd1063,-16'd15,16'd976,-16'd643,-16'd1884,-16'd1858,-16'd3132,-16'd375,-16'd968,-16'd906,16'd270,16'd407,16'd841,-16'd4943,-16'd1836,16'd479,16'd3299,16'd2165,16'd176,-16'd1762,16'd2069,16'd520,16'd2238,-16'd57,-16'd820,16'd563,-16'd589,16'd4407,-16'd416,-16'd1029,-16'd2458,16'd176,-16'd3542,16'd3044,16'd2283,-16'd241,-16'd2033,16'd2617,-16'd1682,16'd227,16'd417,-16'd1230,-16'd947,16'd1708,16'd474,16'd2436,16'd640,-16'd3768,-16'd2612,-16'd153,16'd2472,16'd1515,-16'd1989,-16'd58,-16'd2213,-16'd1958,16'd802,-16'd919,-16'd1596,-16'd2716,16'd4885,-16'd740,16'd1539,16'd858,16'd3201,16'd1980,16'd198,-16'd1960,16'd3012,16'd1645,-16'd3148,-16'd2609,16'd1238,-16'd519,-16'd3026,16'd900,-16'd1682,-16'd1579,-16'd896,-16'd3920,-16'd222,-16'd2210,16'd1021,16'd506,16'd294,16'd341,-16'd234,-16'd384,-16'd1334,16'd3414,16'd2644,16'd2799,16'd893,-16'd1993,-16'd1142,-16'd195,16'd339,16'd710,-16'd1640,16'd634,-16'd1292,-16'd531,16'd2180,16'd963,-16'd519,-16'd3843,-16'd934,-16'd1385,-16'd925,16'd1011,16'd1734,-16'd4736,16'd3566,16'd1478,-16'd3421,16'd993,16'd2049,16'd2302,16'd379,16'd423,16'd1747,16'd6335,-16'd622,16'd1195,-16'd4482,16'd1869,16'd975,-16'd505,16'd2136,-16'd299,16'd4466,-16'd117,16'd108,-16'd2831,-16'd1027,16'd1256,-16'd2833,-16'd671,16'd1492,-16'd112,-16'd3164,16'd789,-16'd2045,-16'd1527,-16'd1794,16'd235,16'd608,-16'd3531,-16'd2910,-16'd690,-16'd2890,16'd3906,16'd1989,-16'd342,-16'd1936,16'd39,16'd2208,16'd512,16'd1200,-16'd147,16'd971,-16'd1058,-16'd5332,-16'd13,-16'd3410,16'd5980,16'd1706,16'd764,-16'd807,16'd2761,16'd210,16'd3218,-16'd486,-16'd737,16'd1342,16'd1969,-16'd678,16'd2382,16'd51,-16'd478,-16'd875,16'd1791,16'd2370,16'd2219,-16'd82,-16'd517,16'd2250,-16'd762,-16'd1459,-16'd2031,16'd2479,16'd2498,-16'd19,-16'd599,16'd1228,-16'd1220,-16'd759,-16'd267,-16'd923,-16'd1444,16'd2785,16'd3216,-16'd4407,16'd817,-16'd724,-16'd3406,-16'd456,-16'd2117,16'd121,16'd338,16'd1014,16'd3844,-16'd2492,16'd606,16'd4502,16'd3870,-16'd423,-16'd1802,16'd3368,-16'd102,-16'd540,-16'd507,-16'd1432,16'd24,-16'd2472,-16'd2227,-16'd1440,16'd1588,-16'd871,16'd9,16'd1166,-16'd2989,-16'd839,16'd1139,16'd1337,-16'd2196,-16'd43,16'd894,16'd3554,16'd1197,16'd1446,16'd426,-16'd5410,-16'd1557,16'd4979,-16'd304,16'd3226,16'd3765,16'd1416,16'd1710,16'd4792,16'd1038,16'd1093,-16'd787,-16'd871,-16'd1799,-16'd571,16'd3459,-16'd1350,16'd2755,-16'd1726,-16'd1639,-16'd82,16'd2885,-16'd2368,-16'd5024,-16'd979,-16'd386,-16'd2659,-16'd1048,-16'd1462,16'd1618,16'd507,16'd2333,-16'd1807,16'd100,-16'd2773,-16'd606,-16'd181,-16'd1174,16'd1617,16'd1626,16'd814,16'd1612,16'd954,16'd185,16'd1294,16'd512,16'd2632,16'd2288,-16'd1201,-16'd1592,-16'd507,-16'd944,-16'd2370,-16'd2136,16'd3976,16'd2732,16'd1072,-16'd2158,16'd620,-16'd2005,-16'd153,16'd2608,-16'd2043,16'd850,16'd1288,16'd479,-16'd2290,16'd520,16'd1235,16'd1637,-16'd1541,-16'd1245,-16'd750,16'd2931,-16'd476,16'd4089,16'd1924,-16'd1052,-16'd1174,16'd1400,16'd3135,-16'd3092,16'd1749,-16'd2604,16'd147,16'd1583,-16'd1789,-16'd4746,16'd1725,-16'd4174,16'd1624,-16'd1426,-16'd316,-16'd1741,16'd2192,-16'd2996,-16'd182,16'd5628,-16'd980,-16'd825,16'd3177,16'd3438,-16'd2510,16'd188,16'd1093,-16'd761,-16'd1153,-16'd3307,16'd718,16'd2320,16'd754,16'd684,16'd4185,-16'd1109,-16'd2234,-16'd51,-16'd2938,-16'd1052,16'd3272,-16'd1553,-16'd4590,-16'd2327,-16'd2893,16'd579,-16'd34,-16'd31,16'd1296,16'd2979,-16'd1727,16'd2145,16'd1099,-16'd1233,16'd1448,16'd3219,16'd3779,-16'd2070,-16'd2842,-16'd1022,-16'd1286,-16'd1519,-16'd1743,-16'd1110,16'd4125,16'd799,-16'd2025,16'd2217,16'd1607,16'd1166,16'd202,-16'd907,-16'd1025,-16'd1899,-16'd1620,-16'd4517,16'd1332,-16'd1556,16'd326,-16'd1421,16'd180,16'd1520,16'd680,-16'd378,-16'd3763,-16'd284,16'd441,-16'd1637,-16'd2576,16'd226,16'd3880,-16'd1068,16'd4440,16'd855,-16'd471,-16'd550,-16'd733,16'd207,-16'd2820,-16'd1741,-16'd2627,-16'd276,-16'd150,16'd888,-16'd573,-16'd710,-16'd3973,16'd2777,-16'd4201,16'd4441,-16'd1350,-16'd2334,16'd1153,16'd2694,16'd2005,16'd953,-16'd98,-16'd1544,-16'd189,-16'd71,16'd123,16'd1751,-16'd1223,16'd2256,16'd307,-16'd2773,16'd1297,16'd1935,-16'd2893,-16'd347,16'd1786,-16'd1473,-16'd34,-16'd1315,-16'd2416,-16'd281,-16'd3480,-16'd865,-16'd44,-16'd296,16'd689,-16'd1588,16'd2744,16'd436,16'd3284,-16'd4387,-16'd1942,16'd444,-16'd2244,16'd1732,-16'd5117,-16'd1724,16'd2229,-16'd2382,16'd721,16'd2100,16'd3307,-16'd745,16'd4641,-16'd980,16'd3292,-16'd3548,-16'd2470,-16'd3169,-16'd4696,16'd1083,16'd890,16'd617,16'd449,-16'd4007,16'd2467,-16'd1836,16'd840,16'd1120,16'd417,16'd1491,16'd258,16'd987,-16'd1643,-16'd2491,-16'd948,-16'd2004,16'd895,-16'd699,16'd415,16'd903,16'd1207,16'd239,-16'd355,-16'd1082,-16'd3368,-16'd141,-16'd998,16'd854,16'd1267,-16'd1073,-16'd2317,16'd953,-16'd475,16'd2805,16'd1915,-16'd214,-16'd3469,16'd505,-16'd1395,-16'd895,-16'd1171,-16'd1870,-16'd2674,-16'd58,-16'd481,16'd3119,-16'd1260,-16'd1593,16'd377,16'd1750,16'd2658,-16'd1048,-16'd647,16'd621,-16'd48,-16'd1163,16'd1360,16'd252,16'd1657,-16'd427,16'd1535,16'd1477,-16'd512,-16'd2684,16'd917,-16'd144,16'd2437,-16'd521,16'd796,-16'd127,-16'd1188,-16'd50,16'd941,-16'd553,-16'd1072,16'd1332,-16'd1853,-16'd2825,16'd227,-16'd2385,-16'd3128,16'd213,16'd1137,-16'd1209,16'd891,-16'd2773,16'd4,-16'd2375,-16'd1933,-16'd1885,-16'd4707,16'd1484,-16'd3571,-16'd62,16'd666,-16'd1879,-16'd74,16'd4434,16'd2079,-16'd885,-16'd1480,-16'd571,-16'd1963,16'd1041,-16'd735,-16'd5068,16'd2791,16'd381,16'd1755,-16'd541,-16'd1079,-16'd1188,-16'd4912,16'd1145,16'd4899,16'd195,16'd1175,16'd2416,16'd628,16'd2187,16'd2784,-16'd2290,16'd1167,16'd2348,16'd113,16'd667,16'd1800,16'd2345,16'd242,16'd1187,-16'd3385,16'd1227,-16'd3205,16'd612,16'd97,-16'd1178,16'd700,16'd1873,16'd419,-16'd1236,-16'd2403,16'd790,-16'd2483,-16'd1852,16'd69,-16'd3866,-16'd314,-16'd3863,16'd3641,16'd332,16'd483,16'd164,16'd2852,16'd89,16'd2431,16'd1722,-16'd4197,-16'd291,-16'd1318,16'd3449,-16'd2651,16'd964,-16'd915,-16'd1902,16'd368,-16'd2918,-16'd1548,16'd3289,-16'd1043,-16'd928,-16'd1135,16'd2728,16'd4229,-16'd2253,-16'd1116,16'd4730,-16'd687,-16'd3720,16'd736,-16'd1851,-16'd4305,16'd267,16'd1083,-16'd2105,-16'd3595,-16'd4294,16'd2703,16'd1297,16'd1995,-16'd2186,16'd1518,-16'd2379,-16'd2137,-16'd644,-16'd175,-16'd2169,16'd919,16'd71,16'd86,16'd3588,-16'd3056,16'd1419,16'd306,-16'd1511,-16'd1891,-16'd3729,-16'd2372,-16'd4226,-16'd608,16'd579,16'd617,-16'd1423,-16'd420,-16'd770,16'd1950,-16'd420,-16'd381,16'd533,16'd721,-16'd7053,-16'd3764,16'd5,16'd1953,-16'd1462,16'd497,-16'd3032,-16'd4605,16'd205,16'd1643,-16'd1398,-16'd432,-16'd941,16'd713,16'd685,-16'd2087,16'd5783,-16'd379,-16'd1031,-16'd1925,16'd1619,-16'd150,16'd64,16'd3449,-16'd693,-16'd1946,-16'd1199,-16'd2596,-16'd3515,16'd1650,16'd2586,16'd713,16'd3808,-16'd3227,-16'd2753,16'd1837,16'd3979,16'd302,16'd349,16'd2377,16'd982,-16'd904,-16'd1274,16'd867,-16'd1068,-16'd2901,16'd361,16'd1030,16'd1198,16'd2682,-16'd567,16'd1107,-16'd2119,16'd5466,16'd988,-16'd986,-16'd1105,16'd1412,-16'd1864,-16'd338,-16'd1297,-16'd253,16'd1852,-16'd264,16'd825,-16'd2469,16'd2650,16'd659,16'd2529,-16'd833,16'd1989,16'd78,16'd2586,16'd967,16'd1335,16'd2927,-16'd352,16'd926,-16'd1277,16'd371,-16'd6350,-16'd1922,16'd299,-16'd2543,-16'd1124,-16'd2198,16'd605,16'd326,16'd635,-16'd170,-16'd2073,-16'd183,-16'd3481,-16'd1403,16'd782,-16'd3248,-16'd321,16'd3881,16'd2328,16'd183,-16'd401,-16'd2156,-16'd103,16'd284,-16'd745,-16'd530,-16'd1451,16'd1223,16'd2084,-16'd3838,16'd551,16'd1313,-16'd2836,16'd45,-16'd1029,16'd62,16'd3042,16'd2037,16'd4377,16'd1968,-16'd381,16'd4212,-16'd1022,-16'd1213,-16'd1555,16'd4042,-16'd178,-16'd872,16'd2730,-16'd3042,16'd1293,-16'd143,-16'd1480,-16'd1787,16'd157,16'd2051,-16'd775,-16'd1826,16'd2230,16'd195,16'd3114,16'd1083,16'd861,16'd81,-16'd475,-16'd260,-16'd3465,-16'd971,-16'd4642,16'd1085,-16'd800,-16'd6361,-16'd1574,16'd2881,16'd4316,-16'd400,16'd1930,-16'd97,16'd2265,-16'd1266,16'd167,-16'd851,16'd1601,16'd233,-16'd961,-16'd1961,-16'd3603,16'd136,16'd2253,16'd4608,16'd1041,-16'd1630,16'd51,16'd1070,-16'd2191,16'd310,-16'd1170,-16'd737,16'd171,-16'd481,-16'd1670,-16'd2406,-16'd1283,-16'd1831,16'd1300,-16'd814,16'd1438,16'd1398,-16'd686,-16'd4188,16'd1632,16'd415,16'd393,16'd4165,-16'd2674,16'd3391,-16'd2111,-16'd2675,-16'd2358,16'd1412,-16'd1798,16'd1531,16'd212,-16'd1646,16'd1510,16'd2041,16'd2808,-16'd3704,-16'd1619,16'd193,-16'd2490,16'd2583,-16'd172,-16'd1007,16'd229,-16'd1338,16'd1443,-16'd1408,-16'd612,16'd1138,-16'd1148,-16'd1950,-16'd746,-16'd1015,-16'd540,16'd494,-16'd1539,16'd1502,16'd1436,-16'd763,16'd677,-16'd360,16'd1097,-16'd742,16'd788,16'd468,16'd1014,-16'd1416,-16'd3044,16'd331,16'd500,-16'd3407,16'd1591,16'd2344,-16'd1083,-16'd1960,-16'd1154,-16'd1963,-16'd1046,16'd422,-16'd147,16'd2561,-16'd1454,-16'd2632,-16'd546,16'd2202,16'd2368,-16'd2791,-16'd1945,16'd2379,16'd1891,-16'd3274,-16'd3692,16'd1891,-16'd814,-16'd2898,16'd17,16'd2098,16'd2902,-16'd4379,16'd2842,16'd36,-16'd1762,16'd586,16'd948,-16'd850,16'd1906,16'd132,16'd2214,16'd2223,16'd249,16'd3529,16'd927,-16'd1324,16'd862,-16'd967,16'd256,-16'd681,16'd336,16'd2852,16'd2937,16'd1925,16'd651,-16'd1777,-16'd264,-16'd457,16'd746,-16'd456,16'd562,16'd2404,16'd3611,16'd1095,-16'd2246,-16'd2245,-16'd466,16'd1190,16'd1069,16'd770,-16'd2381,-16'd2467,16'd2442,16'd34,-16'd200,-16'd2690,16'd1422,16'd71,-16'd345,16'd2684,-16'd1167,-16'd2419,-16'd114,16'd6229,16'd194,-16'd1787,-16'd1485,16'd546,16'd1698,-16'd2484,16'd1196,-16'd704,16'd1588,16'd477,16'd597,16'd2987,16'd118,-16'd3077,16'd3575,16'd747,16'd903,16'd1205,16'd153,-16'd3496,16'd489,-16'd1850,16'd2295,-16'd1847,16'd2884,-16'd531,-16'd3679,16'd44,16'd2898,16'd1226,-16'd1728,16'd1198,-16'd5461,16'd4977,16'd2153,16'd4416,-16'd2989,16'd1072,16'd1856,-16'd1716,-16'd1096,-16'd4273,16'd1546,-16'd2904,16'd2827,16'd572,-16'd2037,16'd1267,-16'd180,16'd843,16'd1937,16'd2022,16'd919,16'd452,16'd2904,16'd3998,16'd1072,16'd4725,-16'd2506,-16'd2832,16'd3106,16'd96,-16'd2384,-16'd344,-16'd761,-16'd705,16'd861,16'd310,-16'd2067,-16'd1430,16'd1186,16'd3974,16'd2230,-16'd1243,-16'd26,16'd983,-16'd2259,-16'd474,-16'd875,16'd724,16'd658,16'd1501,-16'd1244,-16'd298,-16'd1061,16'd779,16'd816,-16'd645,16'd4479,-16'd3273,-16'd3110,-16'd3168,16'd233,-16'd1427,-16'd2412,16'd602,-16'd1959,-16'd1640,16'd4,16'd255,-16'd1467,-16'd2863,-16'd2764,16'd2780,-16'd1428,16'd31,-16'd1594,16'd1622,16'd384,16'd2555,16'd2238,16'd2113,16'd1686,-16'd3106,-16'd854,-16'd998,16'd1888,-16'd317,-16'd1701,16'd1584,-16'd2054,-16'd768,-16'd2613,16'd1549,-16'd709,-16'd1299,-16'd657,-16'd1132,-16'd254,-16'd307,16'd3909,16'd2595,-16'd228,-16'd152,-16'd777,-16'd27,16'd2369,-16'd1625,16'd189,-16'd758,-16'd1002,16'd2212,16'd2275,16'd1461,-16'd1323,16'd1795,16'd175,-16'd124,-16'd809,-16'd2826,-16'd1058,-16'd1046,16'd3127,-16'd5464,-16'd2669,16'd1355,-16'd3992,16'd3551,16'd288,16'd1962,16'd68,16'd3959,-16'd872,-16'd551,16'd554,16'd1749,16'd2790,16'd2205,-16'd1998,16'd1133,-16'd91,-16'd381,16'd1976,16'd31,16'd934,16'd1777,16'd759,-16'd2907,16'd1689,-16'd1062,-16'd502,16'd1115};

*/
    quant Q(
        .snr_idx(4'd10),
        .frac_w(-5'd1),
        .data_in(-16'd2893),
        .llr()
    );
endmodule 
